##
## LEF for PtnCells ;
## created by Encounter v14.28-s033_1 on Thu Jan 19 12:55:16 2017
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fe
  CLASS BLOCK ;
  SIZE 1704.3000 BY 640.8000 ;
  FOREIGN fe 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1701.2100 640.4000 1701.3100 640.8000 ;
    END
  END clk
  PIN rst_async_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 637.6250 1704.3000 637.6750 ;
    END
  END rst_async_n
  PIN i_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1555.8100 0.0000 1555.9100 0.4000 ;
    END
  END i_valid
  PIN i_subsampling
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.2850 640.5800 1701.3350 640.8000 ;
    END
  END i_subsampling
  PIN i_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 637.8250 1704.3000 637.8750 ;
    END
  END i_enable
  PIN i_static_pipe_lat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.2250 1704.3000 638.2750 ;
    END
  END i_static_pipe_lat[9]
  PIN i_static_pipe_lat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.2250 1704.3000 638.2750 ;
    END
  END i_static_pipe_lat[8]
  PIN i_static_pipe_lat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.6850 640.5800 1701.7350 640.8000 ;
    END
  END i_static_pipe_lat[7]
  PIN i_static_pipe_lat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.6850 640.5800 1701.7350 640.8000 ;
    END
  END i_static_pipe_lat[6]
  PIN i_static_pipe_lat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1701.6100 640.4000 1701.7100 640.8000 ;
    END
  END i_static_pipe_lat[5]
  PIN i_static_pipe_lat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.0250 1704.3000 638.0750 ;
    END
  END i_static_pipe_lat[4]
  PIN i_static_pipe_lat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.0250 1704.3000 638.0750 ;
    END
  END i_static_pipe_lat[3]
  PIN i_static_pipe_lat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.4850 640.5800 1701.5350 640.8000 ;
    END
  END i_static_pipe_lat[2]
  PIN i_static_pipe_lat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.4850 640.5800 1701.5350 640.8000 ;
    END
  END i_static_pipe_lat[1]
  PIN i_static_pipe_lat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 637.8250 1704.3000 637.8750 ;
    END
  END i_static_pipe_lat[0]
  PIN i_static_coef[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 640.2250 1704.3000 640.2750 ;
    END
  END i_static_coef[44]
  PIN i_static_coef[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 640.2250 1704.3000 640.2750 ;
    END
  END i_static_coef[43]
  PIN i_static_coef[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 640.0250 1704.3000 640.0750 ;
    END
  END i_static_coef[42]
  PIN i_static_coef[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 640.0250 1704.3000 640.0750 ;
    END
  END i_static_coef[41]
  PIN i_static_coef[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.8250 1704.3000 639.8750 ;
    END
  END i_static_coef[40]
  PIN i_static_coef[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.8250 1704.3000 639.8750 ;
    END
  END i_static_coef[39]
  PIN i_static_coef[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.6250 1704.3000 639.6750 ;
    END
  END i_static_coef[38]
  PIN i_static_coef[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.6250 1704.3000 639.6750 ;
    END
  END i_static_coef[37]
  PIN i_static_coef[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.4250 1704.3000 639.4750 ;
    END
  END i_static_coef[36]
  PIN i_static_coef[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.4250 1704.3000 639.4750 ;
    END
  END i_static_coef[35]
  PIN i_static_coef[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.8850 640.5800 1702.9350 640.8000 ;
    END
  END i_static_coef[34]
  PIN i_static_coef[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.8100 640.4000 1702.9100 640.8000 ;
    END
  END i_static_coef[33]
  PIN i_static_coef[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.2250 1704.3000 639.2750 ;
    END
  END i_static_coef[32]
  PIN i_static_coef[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.2250 1704.3000 639.2750 ;
    END
  END i_static_coef[31]
  PIN i_static_coef[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.6850 640.5800 1702.7350 640.8000 ;
    END
  END i_static_coef[30]
  PIN i_static_coef[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.6850 640.5800 1702.7350 640.8000 ;
    END
  END i_static_coef[29]
  PIN i_static_coef[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.0250 1704.3000 639.0750 ;
    END
  END i_static_coef[28]
  PIN i_static_coef[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.0250 1704.3000 639.0750 ;
    END
  END i_static_coef[27]
  PIN i_static_coef[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.4850 640.5800 1702.5350 640.8000 ;
    END
  END i_static_coef[26]
  PIN i_static_coef[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.4850 640.5800 1702.5350 640.8000 ;
    END
  END i_static_coef[25]
  PIN i_static_coef[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.4100 640.4000 1702.5100 640.8000 ;
    END
  END i_static_coef[24]
  PIN i_static_coef[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.8250 1704.3000 638.8750 ;
    END
  END i_static_coef[23]
  PIN i_static_coef[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.5250 1704.3000 0.5750 ;
    END
  END i_static_coef[22]
  PIN i_static_coef[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.8250 1704.3000 638.8750 ;
    END
  END i_static_coef[21]
  PIN i_static_coef[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.2850 640.5800 1702.3350 640.8000 ;
    END
  END i_static_coef[20]
  PIN i_static_coef[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.5250 1704.3000 0.5750 ;
    END
  END i_static_coef[19]
  PIN i_static_coef[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.6850 0.0000 1703.7350 0.2200 ;
    END
  END i_static_coef[18]
  PIN i_static_coef[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.2850 640.5800 1702.3350 640.8000 ;
    END
  END i_static_coef[17]
  PIN i_static_coef[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.6250 1704.3000 638.6750 ;
    END
  END i_static_coef[16]
  PIN i_static_coef[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.6850 0.0000 1703.7350 0.2200 ;
    END
  END i_static_coef[15]
  PIN i_static_coef[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.6250 1704.3000 638.6750 ;
    END
  END i_static_coef[14]
  PIN i_static_coef[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.7250 1704.3000 0.7750 ;
    END
  END i_static_coef[13]
  PIN i_static_coef[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.7250 1704.3000 0.7750 ;
    END
  END i_static_coef[12]
  PIN i_static_coef[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.4850 0.0000 1703.5350 0.2200 ;
    END
  END i_static_coef[11]
  PIN i_static_coef[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.4850 0.0000 1703.5350 0.2200 ;
    END
  END i_static_coef[10]
  PIN i_static_coef[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.0850 640.5800 1702.1350 640.8000 ;
    END
  END i_static_coef[9]
  PIN i_static_coef[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.9250 1704.3000 0.9750 ;
    END
  END i_static_coef[8]
  PIN i_static_coef[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.9250 1704.3000 0.9750 ;
    END
  END i_static_coef[7]
  PIN i_static_coef[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.0850 640.5800 1702.1350 640.8000 ;
    END
  END i_static_coef[6]
  PIN i_static_coef[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.0100 640.4000 1702.1100 640.8000 ;
    END
  END i_static_coef[5]
  PIN i_static_coef[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.4250 1704.3000 638.4750 ;
    END
  END i_static_coef[4]
  PIN i_static_coef[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.4250 1704.3000 638.4750 ;
    END
  END i_static_coef[3]
  PIN i_static_coef[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.8850 640.5800 1701.9350 640.8000 ;
    END
  END i_static_coef[2]
  PIN i_static_coef[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.8850 640.5800 1701.9350 640.8000 ;
    END
  END i_static_coef[1]
  PIN i_static_coef[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.2850 0.0000 1703.3350 0.2200 ;
    END
  END i_static_coef[0]
  PIN i_data_i[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.9850 0.0000 717.0350 0.2200 ;
    END
  END i_data_i[575]
  PIN i_data_i[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.1850 0.0000 717.2350 0.2200 ;
    END
  END i_data_i[574]
  PIN i_data_i[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.3850 0.0000 717.4350 0.2200 ;
    END
  END i_data_i[573]
  PIN i_data_i[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.5850 0.0000 717.6350 0.2200 ;
    END
  END i_data_i[572]
  PIN i_data_i[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.7850 0.0000 717.8350 0.2200 ;
    END
  END i_data_i[571]
  PIN i_data_i[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.9850 0.0000 718.0350 0.2200 ;
    END
  END i_data_i[570]
  PIN i_data_i[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.3850 0.0000 718.4350 0.2200 ;
    END
  END i_data_i[569]
  PIN i_data_i[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.5850 0.0000 718.6350 0.2200 ;
    END
  END i_data_i[568]
  PIN i_data_i[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.7850 0.0000 718.8350 0.2200 ;
    END
  END i_data_i[567]
  PIN i_data_i[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.9850 0.0000 719.0350 0.2200 ;
    END
  END i_data_i[566]
  PIN i_data_i[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.1850 0.0000 719.2350 0.2200 ;
    END
  END i_data_i[565]
  PIN i_data_i[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.3850 0.0000 719.4350 0.2200 ;
    END
  END i_data_i[564]
  PIN i_data_i[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.5850 0.0000 719.6350 0.2200 ;
    END
  END i_data_i[563]
  PIN i_data_i[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.7850 0.0000 719.8350 0.2200 ;
    END
  END i_data_i[562]
  PIN i_data_i[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.9850 0.0000 720.0350 0.2200 ;
    END
  END i_data_i[561]
  PIN i_data_i[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.1850 0.0000 720.2350 0.2200 ;
    END
  END i_data_i[560]
  PIN i_data_i[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.5850 0.0000 720.6350 0.2200 ;
    END
  END i_data_i[559]
  PIN i_data_i[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.7850 0.0000 720.8350 0.2200 ;
    END
  END i_data_i[558]
  PIN i_data_i[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.9850 0.0000 721.0350 0.2200 ;
    END
  END i_data_i[557]
  PIN i_data_i[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.1850 0.0000 721.2350 0.2200 ;
    END
  END i_data_i[556]
  PIN i_data_i[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.3850 0.0000 721.4350 0.2200 ;
    END
  END i_data_i[555]
  PIN i_data_i[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.5850 0.0000 721.6350 0.2200 ;
    END
  END i_data_i[554]
  PIN i_data_i[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.7850 0.0000 721.8350 0.2200 ;
    END
  END i_data_i[553]
  PIN i_data_i[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.9850 0.0000 722.0350 0.2200 ;
    END
  END i_data_i[552]
  PIN i_data_i[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.1850 0.0000 722.2350 0.2200 ;
    END
  END i_data_i[551]
  PIN i_data_i[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.3850 0.0000 722.4350 0.2200 ;
    END
  END i_data_i[550]
  PIN i_data_i[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.7850 0.0000 722.8350 0.2200 ;
    END
  END i_data_i[549]
  PIN i_data_i[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.9850 0.0000 723.0350 0.2200 ;
    END
  END i_data_i[548]
  PIN i_data_i[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.1850 0.0000 723.2350 0.2200 ;
    END
  END i_data_i[547]
  PIN i_data_i[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.3850 0.0000 723.4350 0.2200 ;
    END
  END i_data_i[546]
  PIN i_data_i[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.5850 0.0000 723.6350 0.2200 ;
    END
  END i_data_i[545]
  PIN i_data_i[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.7850 0.0000 723.8350 0.2200 ;
    END
  END i_data_i[544]
  PIN i_data_i[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.9850 0.0000 724.0350 0.2200 ;
    END
  END i_data_i[543]
  PIN i_data_i[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.1850 0.0000 724.2350 0.2200 ;
    END
  END i_data_i[542]
  PIN i_data_i[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.3850 0.0000 724.4350 0.2200 ;
    END
  END i_data_i[541]
  PIN i_data_i[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.5850 0.0000 724.6350 0.2200 ;
    END
  END i_data_i[540]
  PIN i_data_i[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.9850 0.0000 725.0350 0.2200 ;
    END
  END i_data_i[539]
  PIN i_data_i[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.1850 0.0000 725.2350 0.2200 ;
    END
  END i_data_i[538]
  PIN i_data_i[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.3850 0.0000 725.4350 0.2200 ;
    END
  END i_data_i[537]
  PIN i_data_i[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.5850 0.0000 725.6350 0.2200 ;
    END
  END i_data_i[536]
  PIN i_data_i[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.7850 0.0000 725.8350 0.2200 ;
    END
  END i_data_i[535]
  PIN i_data_i[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.9850 0.0000 726.0350 0.2200 ;
    END
  END i_data_i[534]
  PIN i_data_i[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.1850 0.0000 726.2350 0.2200 ;
    END
  END i_data_i[533]
  PIN i_data_i[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.3850 0.0000 726.4350 0.2200 ;
    END
  END i_data_i[532]
  PIN i_data_i[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.5850 0.0000 726.6350 0.2200 ;
    END
  END i_data_i[531]
  PIN i_data_i[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.7850 0.0000 726.8350 0.2200 ;
    END
  END i_data_i[530]
  PIN i_data_i[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.1850 0.0000 727.2350 0.2200 ;
    END
  END i_data_i[529]
  PIN i_data_i[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.3850 0.0000 727.4350 0.2200 ;
    END
  END i_data_i[528]
  PIN i_data_i[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.5850 0.0000 727.6350 0.2200 ;
    END
  END i_data_i[527]
  PIN i_data_i[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.7850 0.0000 727.8350 0.2200 ;
    END
  END i_data_i[526]
  PIN i_data_i[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.9850 0.0000 728.0350 0.2200 ;
    END
  END i_data_i[525]
  PIN i_data_i[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 728.1850 0.0000 728.2350 0.2200 ;
    END
  END i_data_i[524]
  PIN i_data_i[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.0850 0.0000 732.1350 0.2200 ;
    END
  END i_data_i[523]
  PIN i_data_i[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.2850 0.0000 732.3350 0.2200 ;
    END
  END i_data_i[522]
  PIN i_data_i[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.4850 0.0000 732.5350 0.2200 ;
    END
  END i_data_i[521]
  PIN i_data_i[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.6850 0.0000 732.7350 0.2200 ;
    END
  END i_data_i[520]
  PIN i_data_i[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.0850 0.0000 733.1350 0.2200 ;
    END
  END i_data_i[519]
  PIN i_data_i[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.2850 0.0000 733.3350 0.2200 ;
    END
  END i_data_i[518]
  PIN i_data_i[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.4850 0.0000 733.5350 0.2200 ;
    END
  END i_data_i[517]
  PIN i_data_i[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.6850 0.0000 733.7350 0.2200 ;
    END
  END i_data_i[516]
  PIN i_data_i[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.8850 0.0000 733.9350 0.2200 ;
    END
  END i_data_i[515]
  PIN i_data_i[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.0850 0.0000 734.1350 0.2200 ;
    END
  END i_data_i[514]
  PIN i_data_i[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.2850 0.0000 734.3350 0.2200 ;
    END
  END i_data_i[513]
  PIN i_data_i[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.4850 0.0000 734.5350 0.2200 ;
    END
  END i_data_i[512]
  PIN i_data_i[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.6850 0.0000 734.7350 0.2200 ;
    END
  END i_data_i[511]
  PIN i_data_i[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.8850 0.0000 734.9350 0.2200 ;
    END
  END i_data_i[510]
  PIN i_data_i[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.2850 0.0000 735.3350 0.2200 ;
    END
  END i_data_i[509]
  PIN i_data_i[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.4850 0.0000 735.5350 0.2200 ;
    END
  END i_data_i[508]
  PIN i_data_i[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.6850 0.0000 735.7350 0.2200 ;
    END
  END i_data_i[507]
  PIN i_data_i[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.8850 0.0000 735.9350 0.2200 ;
    END
  END i_data_i[506]
  PIN i_data_i[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.0850 0.0000 736.1350 0.2200 ;
    END
  END i_data_i[505]
  PIN i_data_i[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.2850 0.0000 736.3350 0.2200 ;
    END
  END i_data_i[504]
  PIN i_data_i[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.4850 0.0000 736.5350 0.2200 ;
    END
  END i_data_i[503]
  PIN i_data_i[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.6850 0.0000 736.7350 0.2200 ;
    END
  END i_data_i[502]
  PIN i_data_i[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.8850 0.0000 736.9350 0.2200 ;
    END
  END i_data_i[501]
  PIN i_data_i[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.0850 0.0000 737.1350 0.2200 ;
    END
  END i_data_i[500]
  PIN i_data_i[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.6850 0.0000 737.7350 0.2200 ;
    END
  END i_data_i[499]
  PIN i_data_i[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.8850 0.0000 737.9350 0.2200 ;
    END
  END i_data_i[498]
  PIN i_data_i[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.0850 0.0000 738.1350 0.2200 ;
    END
  END i_data_i[497]
  PIN i_data_i[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.2850 0.0000 738.3350 0.2200 ;
    END
  END i_data_i[496]
  PIN i_data_i[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.4850 0.0000 738.5350 0.2200 ;
    END
  END i_data_i[495]
  PIN i_data_i[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.6850 0.0000 738.7350 0.2200 ;
    END
  END i_data_i[494]
  PIN i_data_i[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.8850 0.0000 738.9350 0.2200 ;
    END
  END i_data_i[493]
  PIN i_data_i[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.0850 0.0000 739.1350 0.2200 ;
    END
  END i_data_i[492]
  PIN i_data_i[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.2850 0.0000 739.3350 0.2200 ;
    END
  END i_data_i[491]
  PIN i_data_i[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.4850 0.0000 739.5350 0.2200 ;
    END
  END i_data_i[490]
  PIN i_data_i[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.8850 0.0000 739.9350 0.2200 ;
    END
  END i_data_i[489]
  PIN i_data_i[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.0850 0.0000 740.1350 0.2200 ;
    END
  END i_data_i[488]
  PIN i_data_i[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.2850 0.0000 740.3350 0.2200 ;
    END
  END i_data_i[487]
  PIN i_data_i[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.4850 0.0000 740.5350 0.2200 ;
    END
  END i_data_i[486]
  PIN i_data_i[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.6850 0.0000 740.7350 0.2200 ;
    END
  END i_data_i[485]
  PIN i_data_i[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.8850 0.0000 740.9350 0.2200 ;
    END
  END i_data_i[484]
  PIN i_data_i[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.0850 0.0000 741.1350 0.2200 ;
    END
  END i_data_i[483]
  PIN i_data_i[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.2850 0.0000 741.3350 0.2200 ;
    END
  END i_data_i[482]
  PIN i_data_i[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.4850 0.0000 741.5350 0.2200 ;
    END
  END i_data_i[481]
  PIN i_data_i[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.6850 0.0000 741.7350 0.2200 ;
    END
  END i_data_i[480]
  PIN i_data_i[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.0850 0.0000 742.1350 0.2200 ;
    END
  END i_data_i[479]
  PIN i_data_i[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.2850 0.0000 742.3350 0.2200 ;
    END
  END i_data_i[478]
  PIN i_data_i[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.4850 0.0000 742.5350 0.2200 ;
    END
  END i_data_i[477]
  PIN i_data_i[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.6850 0.0000 742.7350 0.2200 ;
    END
  END i_data_i[476]
  PIN i_data_i[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.8850 0.0000 742.9350 0.2200 ;
    END
  END i_data_i[475]
  PIN i_data_i[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.0850 0.0000 743.1350 0.2200 ;
    END
  END i_data_i[474]
  PIN i_data_i[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.2850 0.0000 743.3350 0.2200 ;
    END
  END i_data_i[473]
  PIN i_data_i[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.4850 0.0000 743.5350 0.2200 ;
    END
  END i_data_i[472]
  PIN i_data_i[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.6850 0.0000 743.7350 0.2200 ;
    END
  END i_data_i[471]
  PIN i_data_i[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.8850 0.0000 743.9350 0.2200 ;
    END
  END i_data_i[470]
  PIN i_data_i[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.2850 0.0000 744.3350 0.2200 ;
    END
  END i_data_i[469]
  PIN i_data_i[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.4850 0.0000 744.5350 0.2200 ;
    END
  END i_data_i[468]
  PIN i_data_i[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.6850 0.0000 744.7350 0.2200 ;
    END
  END i_data_i[467]
  PIN i_data_i[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.8850 0.0000 744.9350 0.2200 ;
    END
  END i_data_i[466]
  PIN i_data_i[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.0850 0.0000 745.1350 0.2200 ;
    END
  END i_data_i[465]
  PIN i_data_i[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.2850 0.0000 745.3350 0.2200 ;
    END
  END i_data_i[464]
  PIN i_data_i[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.4850 0.0000 745.5350 0.2200 ;
    END
  END i_data_i[463]
  PIN i_data_i[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.6850 0.0000 745.7350 0.2200 ;
    END
  END i_data_i[462]
  PIN i_data_i[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.8850 0.0000 745.9350 0.2200 ;
    END
  END i_data_i[461]
  PIN i_data_i[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.0850 0.0000 746.1350 0.2200 ;
    END
  END i_data_i[460]
  PIN i_data_i[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.4850 0.0000 746.5350 0.2200 ;
    END
  END i_data_i[459]
  PIN i_data_i[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.6850 0.0000 746.7350 0.2200 ;
    END
  END i_data_i[458]
  PIN i_data_i[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.8850 0.0000 746.9350 0.2200 ;
    END
  END i_data_i[457]
  PIN i_data_i[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.0850 0.0000 747.1350 0.2200 ;
    END
  END i_data_i[456]
  PIN i_data_i[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.2850 0.0000 747.3350 0.2200 ;
    END
  END i_data_i[455]
  PIN i_data_i[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.4850 0.0000 747.5350 0.2200 ;
    END
  END i_data_i[454]
  PIN i_data_i[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.6850 0.0000 747.7350 0.2200 ;
    END
  END i_data_i[453]
  PIN i_data_i[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.8850 0.0000 747.9350 0.2200 ;
    END
  END i_data_i[452]
  PIN i_data_i[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.0850 0.0000 748.1350 0.2200 ;
    END
  END i_data_i[451]
  PIN i_data_i[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.2850 0.0000 748.3350 0.2200 ;
    END
  END i_data_i[450]
  PIN i_data_i[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.6850 0.0000 748.7350 0.2200 ;
    END
  END i_data_i[449]
  PIN i_data_i[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.8850 0.0000 748.9350 0.2200 ;
    END
  END i_data_i[448]
  PIN i_data_i[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.0850 0.0000 749.1350 0.2200 ;
    END
  END i_data_i[447]
  PIN i_data_i[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.2850 0.0000 749.3350 0.2200 ;
    END
  END i_data_i[446]
  PIN i_data_i[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.4850 0.0000 749.5350 0.2200 ;
    END
  END i_data_i[445]
  PIN i_data_i[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.6850 0.0000 749.7350 0.2200 ;
    END
  END i_data_i[444]
  PIN i_data_i[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.8850 0.0000 749.9350 0.2200 ;
    END
  END i_data_i[443]
  PIN i_data_i[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.0850 0.0000 750.1350 0.2200 ;
    END
  END i_data_i[442]
  PIN i_data_i[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.2850 0.0000 750.3350 0.2200 ;
    END
  END i_data_i[441]
  PIN i_data_i[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.4850 0.0000 750.5350 0.2200 ;
    END
  END i_data_i[440]
  PIN i_data_i[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.8850 0.0000 750.9350 0.2200 ;
    END
  END i_data_i[439]
  PIN i_data_i[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.0850 0.0000 751.1350 0.2200 ;
    END
  END i_data_i[438]
  PIN i_data_i[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.2850 0.0000 751.3350 0.2200 ;
    END
  END i_data_i[437]
  PIN i_data_i[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.4850 0.0000 751.5350 0.2200 ;
    END
  END i_data_i[436]
  PIN i_data_i[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.6850 0.0000 751.7350 0.2200 ;
    END
  END i_data_i[435]
  PIN i_data_i[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.8850 0.0000 751.9350 0.2200 ;
    END
  END i_data_i[434]
  PIN i_data_i[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.0850 0.0000 752.1350 0.2200 ;
    END
  END i_data_i[433]
  PIN i_data_i[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.2850 0.0000 752.3350 0.2200 ;
    END
  END i_data_i[432]
  PIN i_data_i[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.4850 0.0000 752.5350 0.2200 ;
    END
  END i_data_i[431]
  PIN i_data_i[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.2850 0.0000 756.3350 0.2200 ;
    END
  END i_data_i[430]
  PIN i_data_i[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.6850 0.0000 756.7350 0.2200 ;
    END
  END i_data_i[429]
  PIN i_data_i[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.8850 0.0000 756.9350 0.2200 ;
    END
  END i_data_i[428]
  PIN i_data_i[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.0850 0.0000 757.1350 0.2200 ;
    END
  END i_data_i[427]
  PIN i_data_i[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.2850 0.0000 757.3350 0.2200 ;
    END
  END i_data_i[426]
  PIN i_data_i[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.4850 0.0000 757.5350 0.2200 ;
    END
  END i_data_i[425]
  PIN i_data_i[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.6850 0.0000 757.7350 0.2200 ;
    END
  END i_data_i[424]
  PIN i_data_i[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.8850 0.0000 757.9350 0.2200 ;
    END
  END i_data_i[423]
  PIN i_data_i[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.0850 0.0000 758.1350 0.2200 ;
    END
  END i_data_i[422]
  PIN i_data_i[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.2850 0.0000 758.3350 0.2200 ;
    END
  END i_data_i[421]
  PIN i_data_i[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.4850 0.0000 758.5350 0.2200 ;
    END
  END i_data_i[420]
  PIN i_data_i[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.8850 0.0000 758.9350 0.2200 ;
    END
  END i_data_i[419]
  PIN i_data_i[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.0850 0.0000 759.1350 0.2200 ;
    END
  END i_data_i[418]
  PIN i_data_i[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.2850 0.0000 759.3350 0.2200 ;
    END
  END i_data_i[417]
  PIN i_data_i[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.4850 0.0000 759.5350 0.2200 ;
    END
  END i_data_i[416]
  PIN i_data_i[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.6850 0.0000 759.7350 0.2200 ;
    END
  END i_data_i[415]
  PIN i_data_i[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.8850 0.0000 759.9350 0.2200 ;
    END
  END i_data_i[414]
  PIN i_data_i[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.0850 0.0000 760.1350 0.2200 ;
    END
  END i_data_i[413]
  PIN i_data_i[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.2850 0.0000 760.3350 0.2200 ;
    END
  END i_data_i[412]
  PIN i_data_i[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.4850 0.0000 760.5350 0.2200 ;
    END
  END i_data_i[411]
  PIN i_data_i[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.6850 0.0000 760.7350 0.2200 ;
    END
  END i_data_i[410]
  PIN i_data_i[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.0850 0.0000 761.1350 0.2200 ;
    END
  END i_data_i[409]
  PIN i_data_i[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.2850 0.0000 761.3350 0.2200 ;
    END
  END i_data_i[408]
  PIN i_data_i[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.4850 0.0000 761.5350 0.2200 ;
    END
  END i_data_i[407]
  PIN i_data_i[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.6850 0.0000 761.7350 0.2200 ;
    END
  END i_data_i[406]
  PIN i_data_i[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.8850 0.0000 761.9350 0.2200 ;
    END
  END i_data_i[405]
  PIN i_data_i[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.0850 0.0000 762.1350 0.2200 ;
    END
  END i_data_i[404]
  PIN i_data_i[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.2850 0.0000 762.3350 0.2200 ;
    END
  END i_data_i[403]
  PIN i_data_i[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.4850 0.0000 762.5350 0.2200 ;
    END
  END i_data_i[402]
  PIN i_data_i[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.6850 0.0000 762.7350 0.2200 ;
    END
  END i_data_i[401]
  PIN i_data_i[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.8850 0.0000 762.9350 0.2200 ;
    END
  END i_data_i[400]
  PIN i_data_i[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.4850 0.0000 763.5350 0.2200 ;
    END
  END i_data_i[399]
  PIN i_data_i[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.6850 0.0000 763.7350 0.2200 ;
    END
  END i_data_i[398]
  PIN i_data_i[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.8850 0.0000 763.9350 0.2200 ;
    END
  END i_data_i[397]
  PIN i_data_i[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.0850 0.0000 764.1350 0.2200 ;
    END
  END i_data_i[396]
  PIN i_data_i[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.2850 0.0000 764.3350 0.2200 ;
    END
  END i_data_i[395]
  PIN i_data_i[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.4850 0.0000 764.5350 0.2200 ;
    END
  END i_data_i[394]
  PIN i_data_i[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.6850 0.0000 764.7350 0.2200 ;
    END
  END i_data_i[393]
  PIN i_data_i[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.8850 0.0000 764.9350 0.2200 ;
    END
  END i_data_i[392]
  PIN i_data_i[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.0850 0.0000 765.1350 0.2200 ;
    END
  END i_data_i[391]
  PIN i_data_i[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.2850 0.0000 765.3350 0.2200 ;
    END
  END i_data_i[390]
  PIN i_data_i[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.6850 0.0000 765.7350 0.2200 ;
    END
  END i_data_i[389]
  PIN i_data_i[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.8850 0.0000 765.9350 0.2200 ;
    END
  END i_data_i[388]
  PIN i_data_i[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.0850 0.0000 766.1350 0.2200 ;
    END
  END i_data_i[387]
  PIN i_data_i[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.2850 0.0000 766.3350 0.2200 ;
    END
  END i_data_i[386]
  PIN i_data_i[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.4850 0.0000 766.5350 0.2200 ;
    END
  END i_data_i[385]
  PIN i_data_i[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.6850 0.0000 766.7350 0.2200 ;
    END
  END i_data_i[384]
  PIN i_data_i[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.8850 0.0000 766.9350 0.2200 ;
    END
  END i_data_i[383]
  PIN i_data_i[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.0850 0.0000 767.1350 0.2200 ;
    END
  END i_data_i[382]
  PIN i_data_i[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.2850 0.0000 767.3350 0.2200 ;
    END
  END i_data_i[381]
  PIN i_data_i[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.4850 0.0000 767.5350 0.2200 ;
    END
  END i_data_i[380]
  PIN i_data_i[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.8850 0.0000 767.9350 0.2200 ;
    END
  END i_data_i[379]
  PIN i_data_i[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.0850 0.0000 768.1350 0.2200 ;
    END
  END i_data_i[378]
  PIN i_data_i[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.2850 0.0000 768.3350 0.2200 ;
    END
  END i_data_i[377]
  PIN i_data_i[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.4850 0.0000 768.5350 0.2200 ;
    END
  END i_data_i[376]
  PIN i_data_i[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.6850 0.0000 768.7350 0.2200 ;
    END
  END i_data_i[375]
  PIN i_data_i[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.8850 0.0000 768.9350 0.2200 ;
    END
  END i_data_i[374]
  PIN i_data_i[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.0850 0.0000 769.1350 0.2200 ;
    END
  END i_data_i[373]
  PIN i_data_i[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.2850 0.0000 769.3350 0.2200 ;
    END
  END i_data_i[372]
  PIN i_data_i[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.4850 0.0000 769.5350 0.2200 ;
    END
  END i_data_i[371]
  PIN i_data_i[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.6850 0.0000 769.7350 0.2200 ;
    END
  END i_data_i[370]
  PIN i_data_i[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.0850 0.0000 770.1350 0.2200 ;
    END
  END i_data_i[369]
  PIN i_data_i[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.2850 0.0000 770.3350 0.2200 ;
    END
  END i_data_i[368]
  PIN i_data_i[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.4850 0.0000 770.5350 0.2200 ;
    END
  END i_data_i[367]
  PIN i_data_i[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.6850 0.0000 770.7350 0.2200 ;
    END
  END i_data_i[366]
  PIN i_data_i[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.8850 0.0000 770.9350 0.2200 ;
    END
  END i_data_i[365]
  PIN i_data_i[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.0850 0.0000 771.1350 0.2200 ;
    END
  END i_data_i[364]
  PIN i_data_i[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.2850 0.0000 771.3350 0.2200 ;
    END
  END i_data_i[363]
  PIN i_data_i[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.4850 0.0000 771.5350 0.2200 ;
    END
  END i_data_i[362]
  PIN i_data_i[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.6850 0.0000 771.7350 0.2200 ;
    END
  END i_data_i[361]
  PIN i_data_i[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.8850 0.0000 771.9350 0.2200 ;
    END
  END i_data_i[360]
  PIN i_data_i[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.2850 0.0000 772.3350 0.2200 ;
    END
  END i_data_i[359]
  PIN i_data_i[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.4850 0.0000 772.5350 0.2200 ;
    END
  END i_data_i[358]
  PIN i_data_i[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.6850 0.0000 772.7350 0.2200 ;
    END
  END i_data_i[357]
  PIN i_data_i[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.8850 0.0000 772.9350 0.2200 ;
    END
  END i_data_i[356]
  PIN i_data_i[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.0850 0.0000 773.1350 0.2200 ;
    END
  END i_data_i[355]
  PIN i_data_i[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.2850 0.0000 773.3350 0.2200 ;
    END
  END i_data_i[354]
  PIN i_data_i[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.4850 0.0000 773.5350 0.2200 ;
    END
  END i_data_i[353]
  PIN i_data_i[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.6850 0.0000 773.7350 0.2200 ;
    END
  END i_data_i[352]
  PIN i_data_i[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.8850 0.0000 773.9350 0.2200 ;
    END
  END i_data_i[351]
  PIN i_data_i[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.0850 0.0000 774.1350 0.2200 ;
    END
  END i_data_i[350]
  PIN i_data_i[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.4850 0.0000 774.5350 0.2200 ;
    END
  END i_data_i[349]
  PIN i_data_i[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.6850 0.0000 774.7350 0.2200 ;
    END
  END i_data_i[348]
  PIN i_data_i[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.8850 0.0000 774.9350 0.2200 ;
    END
  END i_data_i[347]
  PIN i_data_i[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.0850 0.0000 775.1350 0.2200 ;
    END
  END i_data_i[346]
  PIN i_data_i[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.2850 0.0000 775.3350 0.2200 ;
    END
  END i_data_i[345]
  PIN i_data_i[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.4850 0.0000 775.5350 0.2200 ;
    END
  END i_data_i[344]
  PIN i_data_i[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.6850 0.0000 775.7350 0.2200 ;
    END
  END i_data_i[343]
  PIN i_data_i[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.8850 0.0000 775.9350 0.2200 ;
    END
  END i_data_i[342]
  PIN i_data_i[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.0850 0.0000 776.1350 0.2200 ;
    END
  END i_data_i[341]
  PIN i_data_i[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.2850 0.0000 776.3350 0.2200 ;
    END
  END i_data_i[340]
  PIN i_data_i[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.6850 0.0000 776.7350 0.2200 ;
    END
  END i_data_i[339]
  PIN i_data_i[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.8850 0.0000 776.9350 0.2200 ;
    END
  END i_data_i[338]
  PIN i_data_i[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.5850 0.0000 780.6350 0.2200 ;
    END
  END i_data_i[337]
  PIN i_data_i[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.7850 0.0000 780.8350 0.2200 ;
    END
  END i_data_i[336]
  PIN i_data_i[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.9850 0.0000 781.0350 0.2200 ;
    END
  END i_data_i[335]
  PIN i_data_i[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.1850 0.0000 781.2350 0.2200 ;
    END
  END i_data_i[334]
  PIN i_data_i[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.3850 0.0000 781.4350 0.2200 ;
    END
  END i_data_i[333]
  PIN i_data_i[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.5850 0.0000 781.6350 0.2200 ;
    END
  END i_data_i[332]
  PIN i_data_i[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.7850 0.0000 781.8350 0.2200 ;
    END
  END i_data_i[331]
  PIN i_data_i[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.9850 0.0000 782.0350 0.2200 ;
    END
  END i_data_i[330]
  PIN i_data_i[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.3850 0.0000 782.4350 0.2200 ;
    END
  END i_data_i[329]
  PIN i_data_i[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.5850 0.0000 782.6350 0.2200 ;
    END
  END i_data_i[328]
  PIN i_data_i[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.7850 0.0000 782.8350 0.2200 ;
    END
  END i_data_i[327]
  PIN i_data_i[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.9850 0.0000 783.0350 0.2200 ;
    END
  END i_data_i[326]
  PIN i_data_i[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.1850 0.0000 783.2350 0.2200 ;
    END
  END i_data_i[325]
  PIN i_data_i[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.3850 0.0000 783.4350 0.2200 ;
    END
  END i_data_i[324]
  PIN i_data_i[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.5850 0.0000 783.6350 0.2200 ;
    END
  END i_data_i[323]
  PIN i_data_i[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.7850 0.0000 783.8350 0.2200 ;
    END
  END i_data_i[322]
  PIN i_data_i[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.9850 0.0000 784.0350 0.2200 ;
    END
  END i_data_i[321]
  PIN i_data_i[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.1850 0.0000 784.2350 0.2200 ;
    END
  END i_data_i[320]
  PIN i_data_i[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.5850 0.0000 784.6350 0.2200 ;
    END
  END i_data_i[319]
  PIN i_data_i[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.7850 0.0000 784.8350 0.2200 ;
    END
  END i_data_i[318]
  PIN i_data_i[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.9850 0.0000 785.0350 0.2200 ;
    END
  END i_data_i[317]
  PIN i_data_i[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.1850 0.0000 785.2350 0.2200 ;
    END
  END i_data_i[316]
  PIN i_data_i[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.3850 0.0000 785.4350 0.2200 ;
    END
  END i_data_i[315]
  PIN i_data_i[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.5850 0.0000 785.6350 0.2200 ;
    END
  END i_data_i[314]
  PIN i_data_i[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.7850 0.0000 785.8350 0.2200 ;
    END
  END i_data_i[313]
  PIN i_data_i[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.9850 0.0000 786.0350 0.2200 ;
    END
  END i_data_i[312]
  PIN i_data_i[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.1850 0.0000 786.2350 0.2200 ;
    END
  END i_data_i[311]
  PIN i_data_i[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.3850 0.0000 786.4350 0.2200 ;
    END
  END i_data_i[310]
  PIN i_data_i[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.7850 0.0000 786.8350 0.2200 ;
    END
  END i_data_i[309]
  PIN i_data_i[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.9850 0.0000 787.0350 0.2200 ;
    END
  END i_data_i[308]
  PIN i_data_i[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.1850 0.0000 787.2350 0.2200 ;
    END
  END i_data_i[307]
  PIN i_data_i[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.3850 0.0000 787.4350 0.2200 ;
    END
  END i_data_i[306]
  PIN i_data_i[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.5850 0.0000 787.6350 0.2200 ;
    END
  END i_data_i[305]
  PIN i_data_i[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.7850 0.0000 787.8350 0.2200 ;
    END
  END i_data_i[304]
  PIN i_data_i[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.9850 0.0000 788.0350 0.2200 ;
    END
  END i_data_i[303]
  PIN i_data_i[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.1850 0.0000 788.2350 0.2200 ;
    END
  END i_data_i[302]
  PIN i_data_i[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.3850 0.0000 788.4350 0.2200 ;
    END
  END i_data_i[301]
  PIN i_data_i[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.5850 0.0000 788.6350 0.2200 ;
    END
  END i_data_i[300]
  PIN i_data_i[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.1850 0.0000 789.2350 0.2200 ;
    END
  END i_data_i[299]
  PIN i_data_i[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.3850 0.0000 789.4350 0.2200 ;
    END
  END i_data_i[298]
  PIN i_data_i[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.5850 0.0000 789.6350 0.2200 ;
    END
  END i_data_i[297]
  PIN i_data_i[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.7850 0.0000 789.8350 0.2200 ;
    END
  END i_data_i[296]
  PIN i_data_i[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.9850 0.0000 790.0350 0.2200 ;
    END
  END i_data_i[295]
  PIN i_data_i[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.1850 0.0000 790.2350 0.2200 ;
    END
  END i_data_i[294]
  PIN i_data_i[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.3850 0.0000 790.4350 0.2200 ;
    END
  END i_data_i[293]
  PIN i_data_i[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.5850 0.0000 790.6350 0.2200 ;
    END
  END i_data_i[292]
  PIN i_data_i[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.7850 0.0000 790.8350 0.2200 ;
    END
  END i_data_i[291]
  PIN i_data_i[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.9850 0.0000 791.0350 0.2200 ;
    END
  END i_data_i[290]
  PIN i_data_i[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.3850 0.0000 791.4350 0.2200 ;
    END
  END i_data_i[289]
  PIN i_data_i[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.5850 0.0000 791.6350 0.2200 ;
    END
  END i_data_i[288]
  PIN i_data_i[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.7850 0.0000 791.8350 0.2200 ;
    END
  END i_data_i[287]
  PIN i_data_i[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.9850 0.0000 792.0350 0.2200 ;
    END
  END i_data_i[286]
  PIN i_data_i[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.1850 0.0000 792.2350 0.2200 ;
    END
  END i_data_i[285]
  PIN i_data_i[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.3850 0.0000 792.4350 0.2200 ;
    END
  END i_data_i[284]
  PIN i_data_i[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.5850 0.0000 792.6350 0.2200 ;
    END
  END i_data_i[283]
  PIN i_data_i[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.7850 0.0000 792.8350 0.2200 ;
    END
  END i_data_i[282]
  PIN i_data_i[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.9850 0.0000 793.0350 0.2200 ;
    END
  END i_data_i[281]
  PIN i_data_i[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.1850 0.0000 793.2350 0.2200 ;
    END
  END i_data_i[280]
  PIN i_data_i[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.5850 0.0000 793.6350 0.2200 ;
    END
  END i_data_i[279]
  PIN i_data_i[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.7850 0.0000 793.8350 0.2200 ;
    END
  END i_data_i[278]
  PIN i_data_i[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.9850 0.0000 794.0350 0.2200 ;
    END
  END i_data_i[277]
  PIN i_data_i[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.1850 0.0000 794.2350 0.2200 ;
    END
  END i_data_i[276]
  PIN i_data_i[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.3850 0.0000 794.4350 0.2200 ;
    END
  END i_data_i[275]
  PIN i_data_i[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.5850 0.0000 794.6350 0.2200 ;
    END
  END i_data_i[274]
  PIN i_data_i[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.7850 0.0000 794.8350 0.2200 ;
    END
  END i_data_i[273]
  PIN i_data_i[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.9850 0.0000 795.0350 0.2200 ;
    END
  END i_data_i[272]
  PIN i_data_i[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.1850 0.0000 795.2350 0.2200 ;
    END
  END i_data_i[271]
  PIN i_data_i[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.3850 0.0000 795.4350 0.2200 ;
    END
  END i_data_i[270]
  PIN i_data_i[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.7850 0.0000 795.8350 0.2200 ;
    END
  END i_data_i[269]
  PIN i_data_i[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.9850 0.0000 796.0350 0.2200 ;
    END
  END i_data_i[268]
  PIN i_data_i[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.1850 0.0000 796.2350 0.2200 ;
    END
  END i_data_i[267]
  PIN i_data_i[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.3850 0.0000 796.4350 0.2200 ;
    END
  END i_data_i[266]
  PIN i_data_i[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.5850 0.0000 796.6350 0.2200 ;
    END
  END i_data_i[265]
  PIN i_data_i[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.7850 0.0000 796.8350 0.2200 ;
    END
  END i_data_i[264]
  PIN i_data_i[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.9850 0.0000 797.0350 0.2200 ;
    END
  END i_data_i[263]
  PIN i_data_i[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.1850 0.0000 797.2350 0.2200 ;
    END
  END i_data_i[262]
  PIN i_data_i[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.3850 0.0000 797.4350 0.2200 ;
    END
  END i_data_i[261]
  PIN i_data_i[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.5850 0.0000 797.6350 0.2200 ;
    END
  END i_data_i[260]
  PIN i_data_i[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.9850 0.0000 798.0350 0.2200 ;
    END
  END i_data_i[259]
  PIN i_data_i[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.1850 0.0000 798.2350 0.2200 ;
    END
  END i_data_i[258]
  PIN i_data_i[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.3850 0.0000 798.4350 0.2200 ;
    END
  END i_data_i[257]
  PIN i_data_i[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.5850 0.0000 798.6350 0.2200 ;
    END
  END i_data_i[256]
  PIN i_data_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.7850 0.0000 798.8350 0.2200 ;
    END
  END i_data_i[255]
  PIN i_data_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.9850 0.0000 799.0350 0.2200 ;
    END
  END i_data_i[254]
  PIN i_data_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.1850 0.0000 799.2350 0.2200 ;
    END
  END i_data_i[253]
  PIN i_data_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.3850 0.0000 799.4350 0.2200 ;
    END
  END i_data_i[252]
  PIN i_data_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.5850 0.0000 799.6350 0.2200 ;
    END
  END i_data_i[251]
  PIN i_data_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.7850 0.0000 799.8350 0.2200 ;
    END
  END i_data_i[250]
  PIN i_data_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.1850 0.0000 800.2350 0.2200 ;
    END
  END i_data_i[249]
  PIN i_data_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.3850 0.0000 800.4350 0.2200 ;
    END
  END i_data_i[248]
  PIN i_data_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.5850 0.0000 800.6350 0.2200 ;
    END
  END i_data_i[247]
  PIN i_data_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.7850 0.0000 800.8350 0.2200 ;
    END
  END i_data_i[246]
  PIN i_data_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.9850 0.0000 801.0350 0.2200 ;
    END
  END i_data_i[245]
  PIN i_data_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 801.1850 0.0000 801.2350 0.2200 ;
    END
  END i_data_i[244]
  PIN i_data_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 804.8850 0.0000 804.9350 0.2200 ;
    END
  END i_data_i[243]
  PIN i_data_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.0850 0.0000 805.1350 0.2200 ;
    END
  END i_data_i[242]
  PIN i_data_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.2850 0.0000 805.3350 0.2200 ;
    END
  END i_data_i[241]
  PIN i_data_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.4850 0.0000 805.5350 0.2200 ;
    END
  END i_data_i[240]
  PIN i_data_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.8850 0.0000 805.9350 0.2200 ;
    END
  END i_data_i[239]
  PIN i_data_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.0850 0.0000 806.1350 0.2200 ;
    END
  END i_data_i[238]
  PIN i_data_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.2850 0.0000 806.3350 0.2200 ;
    END
  END i_data_i[237]
  PIN i_data_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.4850 0.0000 806.5350 0.2200 ;
    END
  END i_data_i[236]
  PIN i_data_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.6850 0.0000 806.7350 0.2200 ;
    END
  END i_data_i[235]
  PIN i_data_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.8850 0.0000 806.9350 0.2200 ;
    END
  END i_data_i[234]
  PIN i_data_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.0850 0.0000 807.1350 0.2200 ;
    END
  END i_data_i[233]
  PIN i_data_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.2850 0.0000 807.3350 0.2200 ;
    END
  END i_data_i[232]
  PIN i_data_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.4850 0.0000 807.5350 0.2200 ;
    END
  END i_data_i[231]
  PIN i_data_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.6850 0.0000 807.7350 0.2200 ;
    END
  END i_data_i[230]
  PIN i_data_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.0850 0.0000 808.1350 0.2200 ;
    END
  END i_data_i[229]
  PIN i_data_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.2850 0.0000 808.3350 0.2200 ;
    END
  END i_data_i[228]
  PIN i_data_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.4850 0.0000 808.5350 0.2200 ;
    END
  END i_data_i[227]
  PIN i_data_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.6850 0.0000 808.7350 0.2200 ;
    END
  END i_data_i[226]
  PIN i_data_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.8850 0.0000 808.9350 0.2200 ;
    END
  END i_data_i[225]
  PIN i_data_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.0850 0.0000 809.1350 0.2200 ;
    END
  END i_data_i[224]
  PIN i_data_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.2850 0.0000 809.3350 0.2200 ;
    END
  END i_data_i[223]
  PIN i_data_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.4850 0.0000 809.5350 0.2200 ;
    END
  END i_data_i[222]
  PIN i_data_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.6850 0.0000 809.7350 0.2200 ;
    END
  END i_data_i[221]
  PIN i_data_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.8850 0.0000 809.9350 0.2200 ;
    END
  END i_data_i[220]
  PIN i_data_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.2850 0.0000 810.3350 0.2200 ;
    END
  END i_data_i[219]
  PIN i_data_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.4850 0.0000 810.5350 0.2200 ;
    END
  END i_data_i[218]
  PIN i_data_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.6850 0.0000 810.7350 0.2200 ;
    END
  END i_data_i[217]
  PIN i_data_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.8850 0.0000 810.9350 0.2200 ;
    END
  END i_data_i[216]
  PIN i_data_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.0850 0.0000 811.1350 0.2200 ;
    END
  END i_data_i[215]
  PIN i_data_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.2850 0.0000 811.3350 0.2200 ;
    END
  END i_data_i[214]
  PIN i_data_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.4850 0.0000 811.5350 0.2200 ;
    END
  END i_data_i[213]
  PIN i_data_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.6850 0.0000 811.7350 0.2200 ;
    END
  END i_data_i[212]
  PIN i_data_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.8850 0.0000 811.9350 0.2200 ;
    END
  END i_data_i[211]
  PIN i_data_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.0850 0.0000 812.1350 0.2200 ;
    END
  END i_data_i[210]
  PIN i_data_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.4850 0.0000 812.5350 0.2200 ;
    END
  END i_data_i[209]
  PIN i_data_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.6850 0.0000 812.7350 0.2200 ;
    END
  END i_data_i[208]
  PIN i_data_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.8850 0.0000 812.9350 0.2200 ;
    END
  END i_data_i[207]
  PIN i_data_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.0850 0.0000 813.1350 0.2200 ;
    END
  END i_data_i[206]
  PIN i_data_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.2850 0.0000 813.3350 0.2200 ;
    END
  END i_data_i[205]
  PIN i_data_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.4850 0.0000 813.5350 0.2200 ;
    END
  END i_data_i[204]
  PIN i_data_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.6850 0.0000 813.7350 0.2200 ;
    END
  END i_data_i[203]
  PIN i_data_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.8850 0.0000 813.9350 0.2200 ;
    END
  END i_data_i[202]
  PIN i_data_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.0850 0.0000 814.1350 0.2200 ;
    END
  END i_data_i[201]
  PIN i_data_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.2850 0.0000 814.3350 0.2200 ;
    END
  END i_data_i[200]
  PIN i_data_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.8850 0.0000 814.9350 0.2200 ;
    END
  END i_data_i[199]
  PIN i_data_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.0850 0.0000 815.1350 0.2200 ;
    END
  END i_data_i[198]
  PIN i_data_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.2850 0.0000 815.3350 0.2200 ;
    END
  END i_data_i[197]
  PIN i_data_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.4850 0.0000 815.5350 0.2200 ;
    END
  END i_data_i[196]
  PIN i_data_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.6850 0.0000 815.7350 0.2200 ;
    END
  END i_data_i[195]
  PIN i_data_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.8850 0.0000 815.9350 0.2200 ;
    END
  END i_data_i[194]
  PIN i_data_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.0850 0.0000 816.1350 0.2200 ;
    END
  END i_data_i[193]
  PIN i_data_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.2850 0.0000 816.3350 0.2200 ;
    END
  END i_data_i[192]
  PIN i_data_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.4850 0.0000 816.5350 0.2200 ;
    END
  END i_data_i[191]
  PIN i_data_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.6850 0.0000 816.7350 0.2200 ;
    END
  END i_data_i[190]
  PIN i_data_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.0850 0.0000 817.1350 0.2200 ;
    END
  END i_data_i[189]
  PIN i_data_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.2850 0.0000 817.3350 0.2200 ;
    END
  END i_data_i[188]
  PIN i_data_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.4850 0.0000 817.5350 0.2200 ;
    END
  END i_data_i[187]
  PIN i_data_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.6850 0.0000 817.7350 0.2200 ;
    END
  END i_data_i[186]
  PIN i_data_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.8850 0.0000 817.9350 0.2200 ;
    END
  END i_data_i[185]
  PIN i_data_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.0850 0.0000 818.1350 0.2200 ;
    END
  END i_data_i[184]
  PIN i_data_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.2850 0.0000 818.3350 0.2200 ;
    END
  END i_data_i[183]
  PIN i_data_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.4850 0.0000 818.5350 0.2200 ;
    END
  END i_data_i[182]
  PIN i_data_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.6850 0.0000 818.7350 0.2200 ;
    END
  END i_data_i[181]
  PIN i_data_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.8850 0.0000 818.9350 0.2200 ;
    END
  END i_data_i[180]
  PIN i_data_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.2850 0.0000 819.3350 0.2200 ;
    END
  END i_data_i[179]
  PIN i_data_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.4850 0.0000 819.5350 0.2200 ;
    END
  END i_data_i[178]
  PIN i_data_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.6850 0.0000 819.7350 0.2200 ;
    END
  END i_data_i[177]
  PIN i_data_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.8850 0.0000 819.9350 0.2200 ;
    END
  END i_data_i[176]
  PIN i_data_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.0850 0.0000 820.1350 0.2200 ;
    END
  END i_data_i[175]
  PIN i_data_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.2850 0.0000 820.3350 0.2200 ;
    END
  END i_data_i[174]
  PIN i_data_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.4850 0.0000 820.5350 0.2200 ;
    END
  END i_data_i[173]
  PIN i_data_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.6850 0.0000 820.7350 0.2200 ;
    END
  END i_data_i[172]
  PIN i_data_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.8850 0.0000 820.9350 0.2200 ;
    END
  END i_data_i[171]
  PIN i_data_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.0850 0.0000 821.1350 0.2200 ;
    END
  END i_data_i[170]
  PIN i_data_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.4850 0.0000 821.5350 0.2200 ;
    END
  END i_data_i[169]
  PIN i_data_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.6850 0.0000 821.7350 0.2200 ;
    END
  END i_data_i[168]
  PIN i_data_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.8850 0.0000 821.9350 0.2200 ;
    END
  END i_data_i[167]
  PIN i_data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.0850 0.0000 822.1350 0.2200 ;
    END
  END i_data_i[166]
  PIN i_data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.2850 0.0000 822.3350 0.2200 ;
    END
  END i_data_i[165]
  PIN i_data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.4850 0.0000 822.5350 0.2200 ;
    END
  END i_data_i[164]
  PIN i_data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.6850 0.0000 822.7350 0.2200 ;
    END
  END i_data_i[163]
  PIN i_data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.8850 0.0000 822.9350 0.2200 ;
    END
  END i_data_i[162]
  PIN i_data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.0850 0.0000 823.1350 0.2200 ;
    END
  END i_data_i[161]
  PIN i_data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.2850 0.0000 823.3350 0.2200 ;
    END
  END i_data_i[160]
  PIN i_data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.6850 0.0000 823.7350 0.2200 ;
    END
  END i_data_i[159]
  PIN i_data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.8850 0.0000 823.9350 0.2200 ;
    END
  END i_data_i[158]
  PIN i_data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.0850 0.0000 824.1350 0.2200 ;
    END
  END i_data_i[157]
  PIN i_data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.2850 0.0000 824.3350 0.2200 ;
    END
  END i_data_i[156]
  PIN i_data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.4850 0.0000 824.5350 0.2200 ;
    END
  END i_data_i[155]
  PIN i_data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.6850 0.0000 824.7350 0.2200 ;
    END
  END i_data_i[154]
  PIN i_data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.8850 0.0000 824.9350 0.2200 ;
    END
  END i_data_i[153]
  PIN i_data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.0850 0.0000 825.1350 0.2200 ;
    END
  END i_data_i[152]
  PIN i_data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.2850 0.0000 825.3350 0.2200 ;
    END
  END i_data_i[151]
  PIN i_data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.4850 0.0000 825.5350 0.2200 ;
    END
  END i_data_i[150]
  PIN i_data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.3850 0.0000 829.4350 0.2200 ;
    END
  END i_data_i[149]
  PIN i_data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.5850 0.0000 829.6350 0.2200 ;
    END
  END i_data_i[148]
  PIN i_data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.7850 0.0000 829.8350 0.2200 ;
    END
  END i_data_i[147]
  PIN i_data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.9850 0.0000 830.0350 0.2200 ;
    END
  END i_data_i[146]
  PIN i_data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.1850 0.0000 830.2350 0.2200 ;
    END
  END i_data_i[145]
  PIN i_data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.3850 0.0000 830.4350 0.2200 ;
    END
  END i_data_i[144]
  PIN i_data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.5850 0.0000 830.6350 0.2200 ;
    END
  END i_data_i[143]
  PIN i_data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.7850 0.0000 830.8350 0.2200 ;
    END
  END i_data_i[142]
  PIN i_data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.9850 0.0000 831.0350 0.2200 ;
    END
  END i_data_i[141]
  PIN i_data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.1850 0.0000 831.2350 0.2200 ;
    END
  END i_data_i[140]
  PIN i_data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.5850 0.0000 831.6350 0.2200 ;
    END
  END i_data_i[139]
  PIN i_data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.7850 0.0000 831.8350 0.2200 ;
    END
  END i_data_i[138]
  PIN i_data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.9850 0.0000 832.0350 0.2200 ;
    END
  END i_data_i[137]
  PIN i_data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.1850 0.0000 832.2350 0.2200 ;
    END
  END i_data_i[136]
  PIN i_data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.3850 0.0000 832.4350 0.2200 ;
    END
  END i_data_i[135]
  PIN i_data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.5850 0.0000 832.6350 0.2200 ;
    END
  END i_data_i[134]
  PIN i_data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.7850 0.0000 832.8350 0.2200 ;
    END
  END i_data_i[133]
  PIN i_data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.9850 0.0000 833.0350 0.2200 ;
    END
  END i_data_i[132]
  PIN i_data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.1850 0.0000 833.2350 0.2200 ;
    END
  END i_data_i[131]
  PIN i_data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.3850 0.0000 833.4350 0.2200 ;
    END
  END i_data_i[130]
  PIN i_data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.7850 0.0000 833.8350 0.2200 ;
    END
  END i_data_i[129]
  PIN i_data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.9850 0.0000 834.0350 0.2200 ;
    END
  END i_data_i[128]
  PIN i_data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.1850 0.0000 834.2350 0.2200 ;
    END
  END i_data_i[127]
  PIN i_data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.3850 0.0000 834.4350 0.2200 ;
    END
  END i_data_i[126]
  PIN i_data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.5850 0.0000 834.6350 0.2200 ;
    END
  END i_data_i[125]
  PIN i_data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.7850 0.0000 834.8350 0.2200 ;
    END
  END i_data_i[124]
  PIN i_data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.9850 0.0000 835.0350 0.2200 ;
    END
  END i_data_i[123]
  PIN i_data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.1850 0.0000 835.2350 0.2200 ;
    END
  END i_data_i[122]
  PIN i_data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.3850 0.0000 835.4350 0.2200 ;
    END
  END i_data_i[121]
  PIN i_data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.5850 0.0000 835.6350 0.2200 ;
    END
  END i_data_i[120]
  PIN i_data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.9850 0.0000 836.0350 0.2200 ;
    END
  END i_data_i[119]
  PIN i_data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.1850 0.0000 836.2350 0.2200 ;
    END
  END i_data_i[118]
  PIN i_data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.3850 0.0000 836.4350 0.2200 ;
    END
  END i_data_i[117]
  PIN i_data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.5850 0.0000 836.6350 0.2200 ;
    END
  END i_data_i[116]
  PIN i_data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.7850 0.0000 836.8350 0.2200 ;
    END
  END i_data_i[115]
  PIN i_data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.9850 0.0000 837.0350 0.2200 ;
    END
  END i_data_i[114]
  PIN i_data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.1850 0.0000 837.2350 0.2200 ;
    END
  END i_data_i[113]
  PIN i_data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.3850 0.0000 837.4350 0.2200 ;
    END
  END i_data_i[112]
  PIN i_data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.5850 0.0000 837.6350 0.2200 ;
    END
  END i_data_i[111]
  PIN i_data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.7850 0.0000 837.8350 0.2200 ;
    END
  END i_data_i[110]
  PIN i_data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.1850 0.0000 838.2350 0.2200 ;
    END
  END i_data_i[109]
  PIN i_data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.3850 0.0000 838.4350 0.2200 ;
    END
  END i_data_i[108]
  PIN i_data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.5850 0.0000 838.6350 0.2200 ;
    END
  END i_data_i[107]
  PIN i_data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.7850 0.0000 838.8350 0.2200 ;
    END
  END i_data_i[106]
  PIN i_data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.9850 0.0000 839.0350 0.2200 ;
    END
  END i_data_i[105]
  PIN i_data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.1850 0.0000 839.2350 0.2200 ;
    END
  END i_data_i[104]
  PIN i_data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.3850 0.0000 839.4350 0.2200 ;
    END
  END i_data_i[103]
  PIN i_data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.5850 0.0000 839.6350 0.2200 ;
    END
  END i_data_i[102]
  PIN i_data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.7850 0.0000 839.8350 0.2200 ;
    END
  END i_data_i[101]
  PIN i_data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.9850 0.0000 840.0350 0.2200 ;
    END
  END i_data_i[100]
  PIN i_data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 703.8850 0.0000 703.9350 0.2200 ;
    END
  END i_data_i[99]
  PIN i_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 707.7850 0.0000 707.8350 0.2200 ;
    END
  END i_data_i[98]
  PIN i_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 707.9850 0.0000 708.0350 0.2200 ;
    END
  END i_data_i[97]
  PIN i_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.1850 0.0000 708.2350 0.2200 ;
    END
  END i_data_i[96]
  PIN i_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.3850 0.0000 708.4350 0.2200 ;
    END
  END i_data_i[95]
  PIN i_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.5850 0.0000 708.6350 0.2200 ;
    END
  END i_data_i[94]
  PIN i_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.7850 0.0000 708.8350 0.2200 ;
    END
  END i_data_i[93]
  PIN i_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.9850 0.0000 709.0350 0.2200 ;
    END
  END i_data_i[92]
  PIN i_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.1850 0.0000 709.2350 0.2200 ;
    END
  END i_data_i[91]
  PIN i_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.3850 0.0000 709.4350 0.2200 ;
    END
  END i_data_i[90]
  PIN i_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.7850 0.0000 709.8350 0.2200 ;
    END
  END i_data_i[89]
  PIN i_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.9850 0.0000 710.0350 0.2200 ;
    END
  END i_data_i[88]
  PIN i_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.1850 0.0000 710.2350 0.2200 ;
    END
  END i_data_i[87]
  PIN i_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.3850 0.0000 710.4350 0.2200 ;
    END
  END i_data_i[86]
  PIN i_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.5850 0.0000 710.6350 0.2200 ;
    END
  END i_data_i[85]
  PIN i_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.7850 0.0000 710.8350 0.2200 ;
    END
  END i_data_i[84]
  PIN i_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.9850 0.0000 711.0350 0.2200 ;
    END
  END i_data_i[83]
  PIN i_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.1850 0.0000 711.2350 0.2200 ;
    END
  END i_data_i[82]
  PIN i_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.3850 0.0000 711.4350 0.2200 ;
    END
  END i_data_i[81]
  PIN i_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.5850 0.0000 711.6350 0.2200 ;
    END
  END i_data_i[80]
  PIN i_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.9850 0.0000 712.0350 0.2200 ;
    END
  END i_data_i[79]
  PIN i_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.1850 0.0000 712.2350 0.2200 ;
    END
  END i_data_i[78]
  PIN i_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.3850 0.0000 712.4350 0.2200 ;
    END
  END i_data_i[77]
  PIN i_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.5850 0.0000 712.6350 0.2200 ;
    END
  END i_data_i[76]
  PIN i_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.7850 0.0000 712.8350 0.2200 ;
    END
  END i_data_i[75]
  PIN i_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.9850 0.0000 713.0350 0.2200 ;
    END
  END i_data_i[74]
  PIN i_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.1850 0.0000 713.2350 0.2200 ;
    END
  END i_data_i[73]
  PIN i_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.3850 0.0000 713.4350 0.2200 ;
    END
  END i_data_i[72]
  PIN i_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.5850 0.0000 713.6350 0.2200 ;
    END
  END i_data_i[71]
  PIN i_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.7850 0.0000 713.8350 0.2200 ;
    END
  END i_data_i[70]
  PIN i_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.1850 0.0000 714.2350 0.2200 ;
    END
  END i_data_i[69]
  PIN i_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.3850 0.0000 714.4350 0.2200 ;
    END
  END i_data_i[68]
  PIN i_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.5850 0.0000 714.6350 0.2200 ;
    END
  END i_data_i[67]
  PIN i_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.7850 0.0000 714.8350 0.2200 ;
    END
  END i_data_i[66]
  PIN i_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.9850 0.0000 715.0350 0.2200 ;
    END
  END i_data_i[65]
  PIN i_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.1850 0.0000 715.2350 0.2200 ;
    END
  END i_data_i[64]
  PIN i_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.3850 0.0000 715.4350 0.2200 ;
    END
  END i_data_i[63]
  PIN i_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.5850 0.0000 715.6350 0.2200 ;
    END
  END i_data_i[62]
  PIN i_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.7850 0.0000 715.8350 0.2200 ;
    END
  END i_data_i[61]
  PIN i_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.9850 0.0000 716.0350 0.2200 ;
    END
  END i_data_i[60]
  PIN i_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.3850 0.0000 716.4350 0.2200 ;
    END
  END i_data_i[59]
  PIN i_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.5850 0.0000 716.6350 0.2200 ;
    END
  END i_data_i[58]
  PIN i_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.7850 0.0000 716.8350 0.2200 ;
    END
  END i_data_i[57]
  PIN i_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.1850 0.0000 718.2350 0.2200 ;
    END
  END i_data_i[56]
  PIN i_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.3850 0.0000 720.4350 0.2200 ;
    END
  END i_data_i[55]
  PIN i_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.5850 0.0000 722.6350 0.2200 ;
    END
  END i_data_i[54]
  PIN i_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.7850 0.0000 724.8350 0.2200 ;
    END
  END i_data_i[53]
  PIN i_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.9850 0.0000 727.0350 0.2200 ;
    END
  END i_data_i[52]
  PIN i_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.8850 0.0000 732.9350 0.2200 ;
    END
  END i_data_i[51]
  PIN i_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.0850 0.0000 735.1350 0.2200 ;
    END
  END i_data_i[50]
  PIN i_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.4850 0.0000 737.5350 0.2200 ;
    END
  END i_data_i[49]
  PIN i_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.6850 0.0000 739.7350 0.2200 ;
    END
  END i_data_i[48]
  PIN i_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.8850 0.0000 741.9350 0.2200 ;
    END
  END i_data_i[47]
  PIN i_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.0850 0.0000 744.1350 0.2200 ;
    END
  END i_data_i[46]
  PIN i_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.2850 0.0000 746.3350 0.2200 ;
    END
  END i_data_i[45]
  PIN i_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.4850 0.0000 748.5350 0.2200 ;
    END
  END i_data_i[44]
  PIN i_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.6850 0.0000 750.7350 0.2200 ;
    END
  END i_data_i[43]
  PIN i_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.4850 0.0000 756.5350 0.2200 ;
    END
  END i_data_i[42]
  PIN i_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.6850 0.0000 758.7350 0.2200 ;
    END
  END i_data_i[41]
  PIN i_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.8850 0.0000 760.9350 0.2200 ;
    END
  END i_data_i[40]
  PIN i_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.2850 0.0000 763.3350 0.2200 ;
    END
  END i_data_i[39]
  PIN i_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.4850 0.0000 765.5350 0.2200 ;
    END
  END i_data_i[38]
  PIN i_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.6850 0.0000 767.7350 0.2200 ;
    END
  END i_data_i[37]
  PIN i_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.8850 0.0000 769.9350 0.2200 ;
    END
  END i_data_i[36]
  PIN i_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.0850 0.0000 772.1350 0.2200 ;
    END
  END i_data_i[35]
  PIN i_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.2850 0.0000 774.3350 0.2200 ;
    END
  END i_data_i[34]
  PIN i_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.4850 0.0000 776.5350 0.2200 ;
    END
  END i_data_i[33]
  PIN i_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.1850 0.0000 782.2350 0.2200 ;
    END
  END i_data_i[32]
  PIN i_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.3850 0.0000 784.4350 0.2200 ;
    END
  END i_data_i[31]
  PIN i_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.5850 0.0000 786.6350 0.2200 ;
    END
  END i_data_i[30]
  PIN i_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.9850 0.0000 789.0350 0.2200 ;
    END
  END i_data_i[29]
  PIN i_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.1850 0.0000 791.2350 0.2200 ;
    END
  END i_data_i[28]
  PIN i_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.3850 0.0000 793.4350 0.2200 ;
    END
  END i_data_i[27]
  PIN i_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.5850 0.0000 795.6350 0.2200 ;
    END
  END i_data_i[26]
  PIN i_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.7850 0.0000 797.8350 0.2200 ;
    END
  END i_data_i[25]
  PIN i_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.9850 0.0000 800.0350 0.2200 ;
    END
  END i_data_i[24]
  PIN i_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.6850 0.0000 805.7350 0.2200 ;
    END
  END i_data_i[23]
  PIN i_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.8850 0.0000 807.9350 0.2200 ;
    END
  END i_data_i[22]
  PIN i_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.0850 0.0000 810.1350 0.2200 ;
    END
  END i_data_i[21]
  PIN i_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.2850 0.0000 812.3350 0.2200 ;
    END
  END i_data_i[20]
  PIN i_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.6850 0.0000 814.7350 0.2200 ;
    END
  END i_data_i[19]
  PIN i_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.8850 0.0000 816.9350 0.2200 ;
    END
  END i_data_i[18]
  PIN i_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.0850 0.0000 819.1350 0.2200 ;
    END
  END i_data_i[17]
  PIN i_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.2850 0.0000 821.3350 0.2200 ;
    END
  END i_data_i[16]
  PIN i_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.4850 0.0000 823.5350 0.2200 ;
    END
  END i_data_i[15]
  PIN i_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.1850 0.0000 829.2350 0.2200 ;
    END
  END i_data_i[14]
  PIN i_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.3850 0.0000 831.4350 0.2200 ;
    END
  END i_data_i[13]
  PIN i_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.5850 0.0000 833.6350 0.2200 ;
    END
  END i_data_i[12]
  PIN i_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.7850 0.0000 835.8350 0.2200 ;
    END
  END i_data_i[11]
  PIN i_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.9850 0.0000 838.0350 0.2200 ;
    END
  END i_data_i[10]
  PIN i_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 703.6850 0.0000 703.7350 0.2200 ;
    END
  END i_data_i[9]
  PIN i_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.5850 0.0000 709.6350 0.2200 ;
    END
  END i_data_i[8]
  PIN i_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.7850 0.0000 711.8350 0.2200 ;
    END
  END i_data_i[7]
  PIN i_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.9850 0.0000 714.0350 0.2200 ;
    END
  END i_data_i[6]
  PIN i_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.1850 0.0000 716.2350 0.2200 ;
    END
  END i_data_i[5]
  PIN i_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.2850 0.0000 737.3350 0.2200 ;
    END
  END i_data_i[4]
  PIN i_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.0850 0.0000 763.1350 0.2200 ;
    END
  END i_data_i[3]
  PIN i_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.7850 0.0000 788.8350 0.2200 ;
    END
  END i_data_i[2]
  PIN i_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.4850 0.0000 814.5350 0.2200 ;
    END
  END i_data_i[1]
  PIN i_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.1850 0.0000 840.2350 0.2200 ;
    END
  END i_data_i[0]
  PIN i_data_q[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.5850 0.0000 963.6350 0.2200 ;
    END
  END i_data_q[575]
  PIN i_data_q[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.3850 0.0000 963.4350 0.2200 ;
    END
  END i_data_q[574]
  PIN i_data_q[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.1850 0.0000 963.2350 0.2200 ;
    END
  END i_data_q[573]
  PIN i_data_q[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.9850 0.0000 963.0350 0.2200 ;
    END
  END i_data_q[572]
  PIN i_data_q[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.7850 0.0000 962.8350 0.2200 ;
    END
  END i_data_q[571]
  PIN i_data_q[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.5850 0.0000 962.6350 0.2200 ;
    END
  END i_data_q[570]
  PIN i_data_q[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.1850 0.0000 962.2350 0.2200 ;
    END
  END i_data_q[569]
  PIN i_data_q[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.9850 0.0000 962.0350 0.2200 ;
    END
  END i_data_q[568]
  PIN i_data_q[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.7850 0.0000 961.8350 0.2200 ;
    END
  END i_data_q[567]
  PIN i_data_q[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.5850 0.0000 961.6350 0.2200 ;
    END
  END i_data_q[566]
  PIN i_data_q[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.3850 0.0000 961.4350 0.2200 ;
    END
  END i_data_q[565]
  PIN i_data_q[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.1850 0.0000 961.2350 0.2200 ;
    END
  END i_data_q[564]
  PIN i_data_q[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.9850 0.0000 961.0350 0.2200 ;
    END
  END i_data_q[563]
  PIN i_data_q[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.7850 0.0000 960.8350 0.2200 ;
    END
  END i_data_q[562]
  PIN i_data_q[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.5850 0.0000 960.6350 0.2200 ;
    END
  END i_data_q[561]
  PIN i_data_q[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.3850 0.0000 960.4350 0.2200 ;
    END
  END i_data_q[560]
  PIN i_data_q[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.9850 0.0000 960.0350 0.2200 ;
    END
  END i_data_q[559]
  PIN i_data_q[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.7850 0.0000 959.8350 0.2200 ;
    END
  END i_data_q[558]
  PIN i_data_q[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.5850 0.0000 959.6350 0.2200 ;
    END
  END i_data_q[557]
  PIN i_data_q[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.3850 0.0000 959.4350 0.2200 ;
    END
  END i_data_q[556]
  PIN i_data_q[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.1850 0.0000 959.2350 0.2200 ;
    END
  END i_data_q[555]
  PIN i_data_q[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.9850 0.0000 959.0350 0.2200 ;
    END
  END i_data_q[554]
  PIN i_data_q[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.7850 0.0000 958.8350 0.2200 ;
    END
  END i_data_q[553]
  PIN i_data_q[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.5850 0.0000 958.6350 0.2200 ;
    END
  END i_data_q[552]
  PIN i_data_q[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.3850 0.0000 958.4350 0.2200 ;
    END
  END i_data_q[551]
  PIN i_data_q[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.1850 0.0000 958.2350 0.2200 ;
    END
  END i_data_q[550]
  PIN i_data_q[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.7850 0.0000 957.8350 0.2200 ;
    END
  END i_data_q[549]
  PIN i_data_q[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.5850 0.0000 957.6350 0.2200 ;
    END
  END i_data_q[548]
  PIN i_data_q[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.3850 0.0000 957.4350 0.2200 ;
    END
  END i_data_q[547]
  PIN i_data_q[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.1850 0.0000 957.2350 0.2200 ;
    END
  END i_data_q[546]
  PIN i_data_q[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.9850 0.0000 957.0350 0.2200 ;
    END
  END i_data_q[545]
  PIN i_data_q[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.7850 0.0000 956.8350 0.2200 ;
    END
  END i_data_q[544]
  PIN i_data_q[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.5850 0.0000 956.6350 0.2200 ;
    END
  END i_data_q[543]
  PIN i_data_q[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.3850 0.0000 956.4350 0.2200 ;
    END
  END i_data_q[542]
  PIN i_data_q[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.1850 0.0000 956.2350 0.2200 ;
    END
  END i_data_q[541]
  PIN i_data_q[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.9850 0.0000 956.0350 0.2200 ;
    END
  END i_data_q[540]
  PIN i_data_q[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.5850 0.0000 955.6350 0.2200 ;
    END
  END i_data_q[539]
  PIN i_data_q[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.3850 0.0000 955.4350 0.2200 ;
    END
  END i_data_q[538]
  PIN i_data_q[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.1850 0.0000 955.2350 0.2200 ;
    END
  END i_data_q[537]
  PIN i_data_q[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.9850 0.0000 955.0350 0.2200 ;
    END
  END i_data_q[536]
  PIN i_data_q[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.7850 0.0000 954.8350 0.2200 ;
    END
  END i_data_q[535]
  PIN i_data_q[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.5850 0.0000 954.6350 0.2200 ;
    END
  END i_data_q[534]
  PIN i_data_q[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.3850 0.0000 954.4350 0.2200 ;
    END
  END i_data_q[533]
  PIN i_data_q[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.1850 0.0000 954.2350 0.2200 ;
    END
  END i_data_q[532]
  PIN i_data_q[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.9850 0.0000 954.0350 0.2200 ;
    END
  END i_data_q[531]
  PIN i_data_q[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.7850 0.0000 953.8350 0.2200 ;
    END
  END i_data_q[530]
  PIN i_data_q[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.3850 0.0000 953.4350 0.2200 ;
    END
  END i_data_q[529]
  PIN i_data_q[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.1850 0.0000 953.2350 0.2200 ;
    END
  END i_data_q[528]
  PIN i_data_q[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.9850 0.0000 953.0350 0.2200 ;
    END
  END i_data_q[527]
  PIN i_data_q[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.7850 0.0000 952.8350 0.2200 ;
    END
  END i_data_q[526]
  PIN i_data_q[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.5850 0.0000 952.6350 0.2200 ;
    END
  END i_data_q[525]
  PIN i_data_q[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.3850 0.0000 952.4350 0.2200 ;
    END
  END i_data_q[524]
  PIN i_data_q[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.1850 0.0000 952.2350 0.2200 ;
    END
  END i_data_q[523]
  PIN i_data_q[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.9850 0.0000 952.0350 0.2200 ;
    END
  END i_data_q[522]
  PIN i_data_q[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.7850 0.0000 951.8350 0.2200 ;
    END
  END i_data_q[521]
  PIN i_data_q[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.5850 0.0000 951.6350 0.2200 ;
    END
  END i_data_q[520]
  PIN i_data_q[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.1850 0.0000 951.2350 0.2200 ;
    END
  END i_data_q[519]
  PIN i_data_q[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.9850 0.0000 951.0350 0.2200 ;
    END
  END i_data_q[518]
  PIN i_data_q[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.7850 0.0000 950.8350 0.2200 ;
    END
  END i_data_q[517]
  PIN i_data_q[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.5850 0.0000 950.6350 0.2200 ;
    END
  END i_data_q[516]
  PIN i_data_q[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.3850 0.0000 950.4350 0.2200 ;
    END
  END i_data_q[515]
  PIN i_data_q[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.1850 0.0000 950.2350 0.2200 ;
    END
  END i_data_q[514]
  PIN i_data_q[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 946.3850 0.0000 946.4350 0.2200 ;
    END
  END i_data_q[513]
  PIN i_data_q[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 946.1850 0.0000 946.2350 0.2200 ;
    END
  END i_data_q[512]
  PIN i_data_q[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.9850 0.0000 946.0350 0.2200 ;
    END
  END i_data_q[511]
  PIN i_data_q[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.7850 0.0000 945.8350 0.2200 ;
    END
  END i_data_q[510]
  PIN i_data_q[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.3850 0.0000 945.4350 0.2200 ;
    END
  END i_data_q[509]
  PIN i_data_q[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.1850 0.0000 945.2350 0.2200 ;
    END
  END i_data_q[508]
  PIN i_data_q[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.9850 0.0000 945.0350 0.2200 ;
    END
  END i_data_q[507]
  PIN i_data_q[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.7850 0.0000 944.8350 0.2200 ;
    END
  END i_data_q[506]
  PIN i_data_q[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.5850 0.0000 944.6350 0.2200 ;
    END
  END i_data_q[505]
  PIN i_data_q[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.3850 0.0000 944.4350 0.2200 ;
    END
  END i_data_q[504]
  PIN i_data_q[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.1850 0.0000 944.2350 0.2200 ;
    END
  END i_data_q[503]
  PIN i_data_q[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.9850 0.0000 944.0350 0.2200 ;
    END
  END i_data_q[502]
  PIN i_data_q[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.7850 0.0000 943.8350 0.2200 ;
    END
  END i_data_q[501]
  PIN i_data_q[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.5850 0.0000 943.6350 0.2200 ;
    END
  END i_data_q[500]
  PIN i_data_q[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.9850 0.0000 943.0350 0.2200 ;
    END
  END i_data_q[499]
  PIN i_data_q[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.7850 0.0000 942.8350 0.2200 ;
    END
  END i_data_q[498]
  PIN i_data_q[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.5850 0.0000 942.6350 0.2200 ;
    END
  END i_data_q[497]
  PIN i_data_q[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.3850 0.0000 942.4350 0.2200 ;
    END
  END i_data_q[496]
  PIN i_data_q[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.1850 0.0000 942.2350 0.2200 ;
    END
  END i_data_q[495]
  PIN i_data_q[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.9850 0.0000 942.0350 0.2200 ;
    END
  END i_data_q[494]
  PIN i_data_q[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.7850 0.0000 941.8350 0.2200 ;
    END
  END i_data_q[493]
  PIN i_data_q[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.5850 0.0000 941.6350 0.2200 ;
    END
  END i_data_q[492]
  PIN i_data_q[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.3850 0.0000 941.4350 0.2200 ;
    END
  END i_data_q[491]
  PIN i_data_q[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.1850 0.0000 941.2350 0.2200 ;
    END
  END i_data_q[490]
  PIN i_data_q[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.7850 0.0000 940.8350 0.2200 ;
    END
  END i_data_q[489]
  PIN i_data_q[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.5850 0.0000 940.6350 0.2200 ;
    END
  END i_data_q[488]
  PIN i_data_q[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.3850 0.0000 940.4350 0.2200 ;
    END
  END i_data_q[487]
  PIN i_data_q[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.1850 0.0000 940.2350 0.2200 ;
    END
  END i_data_q[486]
  PIN i_data_q[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.9850 0.0000 940.0350 0.2200 ;
    END
  END i_data_q[485]
  PIN i_data_q[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.7850 0.0000 939.8350 0.2200 ;
    END
  END i_data_q[484]
  PIN i_data_q[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.5850 0.0000 939.6350 0.2200 ;
    END
  END i_data_q[483]
  PIN i_data_q[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.3850 0.0000 939.4350 0.2200 ;
    END
  END i_data_q[482]
  PIN i_data_q[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.1850 0.0000 939.2350 0.2200 ;
    END
  END i_data_q[481]
  PIN i_data_q[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.9850 0.0000 939.0350 0.2200 ;
    END
  END i_data_q[480]
  PIN i_data_q[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.5850 0.0000 938.6350 0.2200 ;
    END
  END i_data_q[479]
  PIN i_data_q[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.3850 0.0000 938.4350 0.2200 ;
    END
  END i_data_q[478]
  PIN i_data_q[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.1850 0.0000 938.2350 0.2200 ;
    END
  END i_data_q[477]
  PIN i_data_q[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.9850 0.0000 938.0350 0.2200 ;
    END
  END i_data_q[476]
  PIN i_data_q[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.7850 0.0000 937.8350 0.2200 ;
    END
  END i_data_q[475]
  PIN i_data_q[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.5850 0.0000 937.6350 0.2200 ;
    END
  END i_data_q[474]
  PIN i_data_q[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.3850 0.0000 937.4350 0.2200 ;
    END
  END i_data_q[473]
  PIN i_data_q[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.1850 0.0000 937.2350 0.2200 ;
    END
  END i_data_q[472]
  PIN i_data_q[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.9850 0.0000 937.0350 0.2200 ;
    END
  END i_data_q[471]
  PIN i_data_q[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.7850 0.0000 936.8350 0.2200 ;
    END
  END i_data_q[470]
  PIN i_data_q[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.3850 0.0000 936.4350 0.2200 ;
    END
  END i_data_q[469]
  PIN i_data_q[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.1850 0.0000 936.2350 0.2200 ;
    END
  END i_data_q[468]
  PIN i_data_q[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.9850 0.0000 936.0350 0.2200 ;
    END
  END i_data_q[467]
  PIN i_data_q[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.7850 0.0000 935.8350 0.2200 ;
    END
  END i_data_q[466]
  PIN i_data_q[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.5850 0.0000 935.6350 0.2200 ;
    END
  END i_data_q[465]
  PIN i_data_q[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.3850 0.0000 935.4350 0.2200 ;
    END
  END i_data_q[464]
  PIN i_data_q[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.1850 0.0000 935.2350 0.2200 ;
    END
  END i_data_q[463]
  PIN i_data_q[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.9850 0.0000 935.0350 0.2200 ;
    END
  END i_data_q[462]
  PIN i_data_q[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.7850 0.0000 934.8350 0.2200 ;
    END
  END i_data_q[461]
  PIN i_data_q[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.5850 0.0000 934.6350 0.2200 ;
    END
  END i_data_q[460]
  PIN i_data_q[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.1850 0.0000 934.2350 0.2200 ;
    END
  END i_data_q[459]
  PIN i_data_q[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.9850 0.0000 934.0350 0.2200 ;
    END
  END i_data_q[458]
  PIN i_data_q[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.7850 0.0000 933.8350 0.2200 ;
    END
  END i_data_q[457]
  PIN i_data_q[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.5850 0.0000 933.6350 0.2200 ;
    END
  END i_data_q[456]
  PIN i_data_q[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.3850 0.0000 933.4350 0.2200 ;
    END
  END i_data_q[455]
  PIN i_data_q[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.1850 0.0000 933.2350 0.2200 ;
    END
  END i_data_q[454]
  PIN i_data_q[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.9850 0.0000 933.0350 0.2200 ;
    END
  END i_data_q[453]
  PIN i_data_q[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.7850 0.0000 932.8350 0.2200 ;
    END
  END i_data_q[452]
  PIN i_data_q[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.5850 0.0000 932.6350 0.2200 ;
    END
  END i_data_q[451]
  PIN i_data_q[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.3850 0.0000 932.4350 0.2200 ;
    END
  END i_data_q[450]
  PIN i_data_q[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.9850 0.0000 932.0350 0.2200 ;
    END
  END i_data_q[449]
  PIN i_data_q[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.7850 0.0000 931.8350 0.2200 ;
    END
  END i_data_q[448]
  PIN i_data_q[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.5850 0.0000 931.6350 0.2200 ;
    END
  END i_data_q[447]
  PIN i_data_q[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.3850 0.0000 931.4350 0.2200 ;
    END
  END i_data_q[446]
  PIN i_data_q[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.1850 0.0000 931.2350 0.2200 ;
    END
  END i_data_q[445]
  PIN i_data_q[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.9850 0.0000 931.0350 0.2200 ;
    END
  END i_data_q[444]
  PIN i_data_q[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.7850 0.0000 930.8350 0.2200 ;
    END
  END i_data_q[443]
  PIN i_data_q[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.5850 0.0000 930.6350 0.2200 ;
    END
  END i_data_q[442]
  PIN i_data_q[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.3850 0.0000 930.4350 0.2200 ;
    END
  END i_data_q[441]
  PIN i_data_q[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.1850 0.0000 930.2350 0.2200 ;
    END
  END i_data_q[440]
  PIN i_data_q[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.7850 0.0000 929.8350 0.2200 ;
    END
  END i_data_q[439]
  PIN i_data_q[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.5850 0.0000 929.6350 0.2200 ;
    END
  END i_data_q[438]
  PIN i_data_q[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.3850 0.0000 929.4350 0.2200 ;
    END
  END i_data_q[437]
  PIN i_data_q[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.1850 0.0000 929.2350 0.2200 ;
    END
  END i_data_q[436]
  PIN i_data_q[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.9850 0.0000 929.0350 0.2200 ;
    END
  END i_data_q[435]
  PIN i_data_q[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.7850 0.0000 928.8350 0.2200 ;
    END
  END i_data_q[434]
  PIN i_data_q[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.5850 0.0000 928.6350 0.2200 ;
    END
  END i_data_q[433]
  PIN i_data_q[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.3850 0.0000 928.4350 0.2200 ;
    END
  END i_data_q[432]
  PIN i_data_q[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.1850 0.0000 928.2350 0.2200 ;
    END
  END i_data_q[431]
  PIN i_data_q[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.9850 0.0000 928.0350 0.2200 ;
    END
  END i_data_q[430]
  PIN i_data_q[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.5850 0.0000 927.6350 0.2200 ;
    END
  END i_data_q[429]
  PIN i_data_q[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.3850 0.0000 927.4350 0.2200 ;
    END
  END i_data_q[428]
  PIN i_data_q[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.1850 0.0000 927.2350 0.2200 ;
    END
  END i_data_q[427]
  PIN i_data_q[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.9850 0.0000 927.0350 0.2200 ;
    END
  END i_data_q[426]
  PIN i_data_q[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.7850 0.0000 926.8350 0.2200 ;
    END
  END i_data_q[425]
  PIN i_data_q[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.5850 0.0000 926.6350 0.2200 ;
    END
  END i_data_q[424]
  PIN i_data_q[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.3850 0.0000 926.4350 0.2200 ;
    END
  END i_data_q[423]
  PIN i_data_q[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.1850 0.0000 926.2350 0.2200 ;
    END
  END i_data_q[422]
  PIN i_data_q[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 922.3850 0.0000 922.4350 0.2200 ;
    END
  END i_data_q[421]
  PIN i_data_q[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 922.1850 0.0000 922.2350 0.2200 ;
    END
  END i_data_q[420]
  PIN i_data_q[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.7850 0.0000 921.8350 0.2200 ;
    END
  END i_data_q[419]
  PIN i_data_q[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.5850 0.0000 921.6350 0.2200 ;
    END
  END i_data_q[418]
  PIN i_data_q[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.3850 0.0000 921.4350 0.2200 ;
    END
  END i_data_q[417]
  PIN i_data_q[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.1850 0.0000 921.2350 0.2200 ;
    END
  END i_data_q[416]
  PIN i_data_q[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.9850 0.0000 921.0350 0.2200 ;
    END
  END i_data_q[415]
  PIN i_data_q[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.7850 0.0000 920.8350 0.2200 ;
    END
  END i_data_q[414]
  PIN i_data_q[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.5850 0.0000 920.6350 0.2200 ;
    END
  END i_data_q[413]
  PIN i_data_q[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.3850 0.0000 920.4350 0.2200 ;
    END
  END i_data_q[412]
  PIN i_data_q[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.1850 0.0000 920.2350 0.2200 ;
    END
  END i_data_q[411]
  PIN i_data_q[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.9850 0.0000 920.0350 0.2200 ;
    END
  END i_data_q[410]
  PIN i_data_q[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.5850 0.0000 919.6350 0.2200 ;
    END
  END i_data_q[409]
  PIN i_data_q[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.3850 0.0000 919.4350 0.2200 ;
    END
  END i_data_q[408]
  PIN i_data_q[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.1850 0.0000 919.2350 0.2200 ;
    END
  END i_data_q[407]
  PIN i_data_q[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.9850 0.0000 919.0350 0.2200 ;
    END
  END i_data_q[406]
  PIN i_data_q[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.7850 0.0000 918.8350 0.2200 ;
    END
  END i_data_q[405]
  PIN i_data_q[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.5850 0.0000 918.6350 0.2200 ;
    END
  END i_data_q[404]
  PIN i_data_q[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.3850 0.0000 918.4350 0.2200 ;
    END
  END i_data_q[403]
  PIN i_data_q[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.1850 0.0000 918.2350 0.2200 ;
    END
  END i_data_q[402]
  PIN i_data_q[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.9850 0.0000 918.0350 0.2200 ;
    END
  END i_data_q[401]
  PIN i_data_q[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.7850 0.0000 917.8350 0.2200 ;
    END
  END i_data_q[400]
  PIN i_data_q[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.1850 0.0000 917.2350 0.2200 ;
    END
  END i_data_q[399]
  PIN i_data_q[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.9850 0.0000 917.0350 0.2200 ;
    END
  END i_data_q[398]
  PIN i_data_q[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.7850 0.0000 916.8350 0.2200 ;
    END
  END i_data_q[397]
  PIN i_data_q[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.5850 0.0000 916.6350 0.2200 ;
    END
  END i_data_q[396]
  PIN i_data_q[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.3850 0.0000 916.4350 0.2200 ;
    END
  END i_data_q[395]
  PIN i_data_q[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.1850 0.0000 916.2350 0.2200 ;
    END
  END i_data_q[394]
  PIN i_data_q[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.9850 0.0000 916.0350 0.2200 ;
    END
  END i_data_q[393]
  PIN i_data_q[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.7850 0.0000 915.8350 0.2200 ;
    END
  END i_data_q[392]
  PIN i_data_q[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.5850 0.0000 915.6350 0.2200 ;
    END
  END i_data_q[391]
  PIN i_data_q[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.3850 0.0000 915.4350 0.2200 ;
    END
  END i_data_q[390]
  PIN i_data_q[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.9850 0.0000 915.0350 0.2200 ;
    END
  END i_data_q[389]
  PIN i_data_q[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.7850 0.0000 914.8350 0.2200 ;
    END
  END i_data_q[388]
  PIN i_data_q[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.5850 0.0000 914.6350 0.2200 ;
    END
  END i_data_q[387]
  PIN i_data_q[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.3850 0.0000 914.4350 0.2200 ;
    END
  END i_data_q[386]
  PIN i_data_q[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.1850 0.0000 914.2350 0.2200 ;
    END
  END i_data_q[385]
  PIN i_data_q[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.9850 0.0000 914.0350 0.2200 ;
    END
  END i_data_q[384]
  PIN i_data_q[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.7850 0.0000 913.8350 0.2200 ;
    END
  END i_data_q[383]
  PIN i_data_q[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.5850 0.0000 913.6350 0.2200 ;
    END
  END i_data_q[382]
  PIN i_data_q[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.3850 0.0000 913.4350 0.2200 ;
    END
  END i_data_q[381]
  PIN i_data_q[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.1850 0.0000 913.2350 0.2200 ;
    END
  END i_data_q[380]
  PIN i_data_q[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.7850 0.0000 912.8350 0.2200 ;
    END
  END i_data_q[379]
  PIN i_data_q[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.5850 0.0000 912.6350 0.2200 ;
    END
  END i_data_q[378]
  PIN i_data_q[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.3850 0.0000 912.4350 0.2200 ;
    END
  END i_data_q[377]
  PIN i_data_q[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.1850 0.0000 912.2350 0.2200 ;
    END
  END i_data_q[376]
  PIN i_data_q[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.9850 0.0000 912.0350 0.2200 ;
    END
  END i_data_q[375]
  PIN i_data_q[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.7850 0.0000 911.8350 0.2200 ;
    END
  END i_data_q[374]
  PIN i_data_q[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.5850 0.0000 911.6350 0.2200 ;
    END
  END i_data_q[373]
  PIN i_data_q[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.3850 0.0000 911.4350 0.2200 ;
    END
  END i_data_q[372]
  PIN i_data_q[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.1850 0.0000 911.2350 0.2200 ;
    END
  END i_data_q[371]
  PIN i_data_q[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.9850 0.0000 911.0350 0.2200 ;
    END
  END i_data_q[370]
  PIN i_data_q[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.5850 0.0000 910.6350 0.2200 ;
    END
  END i_data_q[369]
  PIN i_data_q[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.3850 0.0000 910.4350 0.2200 ;
    END
  END i_data_q[368]
  PIN i_data_q[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.1850 0.0000 910.2350 0.2200 ;
    END
  END i_data_q[367]
  PIN i_data_q[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.9850 0.0000 910.0350 0.2200 ;
    END
  END i_data_q[366]
  PIN i_data_q[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.7850 0.0000 909.8350 0.2200 ;
    END
  END i_data_q[365]
  PIN i_data_q[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.5850 0.0000 909.6350 0.2200 ;
    END
  END i_data_q[364]
  PIN i_data_q[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.3850 0.0000 909.4350 0.2200 ;
    END
  END i_data_q[363]
  PIN i_data_q[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.1850 0.0000 909.2350 0.2200 ;
    END
  END i_data_q[362]
  PIN i_data_q[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.9850 0.0000 909.0350 0.2200 ;
    END
  END i_data_q[361]
  PIN i_data_q[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.7850 0.0000 908.8350 0.2200 ;
    END
  END i_data_q[360]
  PIN i_data_q[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.3850 0.0000 908.4350 0.2200 ;
    END
  END i_data_q[359]
  PIN i_data_q[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.1850 0.0000 908.2350 0.2200 ;
    END
  END i_data_q[358]
  PIN i_data_q[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.9850 0.0000 908.0350 0.2200 ;
    END
  END i_data_q[357]
  PIN i_data_q[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.7850 0.0000 907.8350 0.2200 ;
    END
  END i_data_q[356]
  PIN i_data_q[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.5850 0.0000 907.6350 0.2200 ;
    END
  END i_data_q[355]
  PIN i_data_q[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.3850 0.0000 907.4350 0.2200 ;
    END
  END i_data_q[354]
  PIN i_data_q[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.1850 0.0000 907.2350 0.2200 ;
    END
  END i_data_q[353]
  PIN i_data_q[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.9850 0.0000 907.0350 0.2200 ;
    END
  END i_data_q[352]
  PIN i_data_q[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.7850 0.0000 906.8350 0.2200 ;
    END
  END i_data_q[351]
  PIN i_data_q[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.5850 0.0000 906.6350 0.2200 ;
    END
  END i_data_q[350]
  PIN i_data_q[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.1850 0.0000 906.2350 0.2200 ;
    END
  END i_data_q[349]
  PIN i_data_q[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.9850 0.0000 906.0350 0.2200 ;
    END
  END i_data_q[348]
  PIN i_data_q[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.7850 0.0000 905.8350 0.2200 ;
    END
  END i_data_q[347]
  PIN i_data_q[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.5850 0.0000 905.6350 0.2200 ;
    END
  END i_data_q[346]
  PIN i_data_q[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.3850 0.0000 905.4350 0.2200 ;
    END
  END i_data_q[345]
  PIN i_data_q[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.1850 0.0000 905.2350 0.2200 ;
    END
  END i_data_q[344]
  PIN i_data_q[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.9850 0.0000 905.0350 0.2200 ;
    END
  END i_data_q[343]
  PIN i_data_q[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.7850 0.0000 904.8350 0.2200 ;
    END
  END i_data_q[342]
  PIN i_data_q[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.5850 0.0000 904.6350 0.2200 ;
    END
  END i_data_q[341]
  PIN i_data_q[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.3850 0.0000 904.4350 0.2200 ;
    END
  END i_data_q[340]
  PIN i_data_q[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.9850 0.0000 904.0350 0.2200 ;
    END
  END i_data_q[339]
  PIN i_data_q[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.7850 0.0000 903.8350 0.2200 ;
    END
  END i_data_q[338]
  PIN i_data_q[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.5850 0.0000 903.6350 0.2200 ;
    END
  END i_data_q[337]
  PIN i_data_q[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.3850 0.0000 903.4350 0.2200 ;
    END
  END i_data_q[336]
  PIN i_data_q[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.1850 0.0000 903.2350 0.2200 ;
    END
  END i_data_q[335]
  PIN i_data_q[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.9850 0.0000 903.0350 0.2200 ;
    END
  END i_data_q[334]
  PIN i_data_q[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.7850 0.0000 902.8350 0.2200 ;
    END
  END i_data_q[333]
  PIN i_data_q[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.5850 0.0000 902.6350 0.2200 ;
    END
  END i_data_q[332]
  PIN i_data_q[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.3850 0.0000 902.4350 0.2200 ;
    END
  END i_data_q[331]
  PIN i_data_q[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.1850 0.0000 902.2350 0.2200 ;
    END
  END i_data_q[330]
  PIN i_data_q[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 898.1850 0.0000 898.2350 0.2200 ;
    END
  END i_data_q[329]
  PIN i_data_q[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.9850 0.0000 898.0350 0.2200 ;
    END
  END i_data_q[328]
  PIN i_data_q[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.7850 0.0000 897.8350 0.2200 ;
    END
  END i_data_q[327]
  PIN i_data_q[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.5850 0.0000 897.6350 0.2200 ;
    END
  END i_data_q[326]
  PIN i_data_q[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.3850 0.0000 897.4350 0.2200 ;
    END
  END i_data_q[325]
  PIN i_data_q[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.1850 0.0000 897.2350 0.2200 ;
    END
  END i_data_q[324]
  PIN i_data_q[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.9850 0.0000 897.0350 0.2200 ;
    END
  END i_data_q[323]
  PIN i_data_q[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.7850 0.0000 896.8350 0.2200 ;
    END
  END i_data_q[322]
  PIN i_data_q[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.5850 0.0000 896.6350 0.2200 ;
    END
  END i_data_q[321]
  PIN i_data_q[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.3850 0.0000 896.4350 0.2200 ;
    END
  END i_data_q[320]
  PIN i_data_q[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.9850 0.0000 896.0350 0.2200 ;
    END
  END i_data_q[319]
  PIN i_data_q[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.7850 0.0000 895.8350 0.2200 ;
    END
  END i_data_q[318]
  PIN i_data_q[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.5850 0.0000 895.6350 0.2200 ;
    END
  END i_data_q[317]
  PIN i_data_q[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.3850 0.0000 895.4350 0.2200 ;
    END
  END i_data_q[316]
  PIN i_data_q[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.1850 0.0000 895.2350 0.2200 ;
    END
  END i_data_q[315]
  PIN i_data_q[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.9850 0.0000 895.0350 0.2200 ;
    END
  END i_data_q[314]
  PIN i_data_q[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.7850 0.0000 894.8350 0.2200 ;
    END
  END i_data_q[313]
  PIN i_data_q[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.5850 0.0000 894.6350 0.2200 ;
    END
  END i_data_q[312]
  PIN i_data_q[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.3850 0.0000 894.4350 0.2200 ;
    END
  END i_data_q[311]
  PIN i_data_q[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.1850 0.0000 894.2350 0.2200 ;
    END
  END i_data_q[310]
  PIN i_data_q[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.7850 0.0000 893.8350 0.2200 ;
    END
  END i_data_q[309]
  PIN i_data_q[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.5850 0.0000 893.6350 0.2200 ;
    END
  END i_data_q[308]
  PIN i_data_q[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.3850 0.0000 893.4350 0.2200 ;
    END
  END i_data_q[307]
  PIN i_data_q[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.1850 0.0000 893.2350 0.2200 ;
    END
  END i_data_q[306]
  PIN i_data_q[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.9850 0.0000 893.0350 0.2200 ;
    END
  END i_data_q[305]
  PIN i_data_q[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.7850 0.0000 892.8350 0.2200 ;
    END
  END i_data_q[304]
  PIN i_data_q[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.5850 0.0000 892.6350 0.2200 ;
    END
  END i_data_q[303]
  PIN i_data_q[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.3850 0.0000 892.4350 0.2200 ;
    END
  END i_data_q[302]
  PIN i_data_q[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.1850 0.0000 892.2350 0.2200 ;
    END
  END i_data_q[301]
  PIN i_data_q[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.9850 0.0000 892.0350 0.2200 ;
    END
  END i_data_q[300]
  PIN i_data_q[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.3850 0.0000 891.4350 0.2200 ;
    END
  END i_data_q[299]
  PIN i_data_q[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.1850 0.0000 891.2350 0.2200 ;
    END
  END i_data_q[298]
  PIN i_data_q[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.9850 0.0000 891.0350 0.2200 ;
    END
  END i_data_q[297]
  PIN i_data_q[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.7850 0.0000 890.8350 0.2200 ;
    END
  END i_data_q[296]
  PIN i_data_q[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.5850 0.0000 890.6350 0.2200 ;
    END
  END i_data_q[295]
  PIN i_data_q[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.3850 0.0000 890.4350 0.2200 ;
    END
  END i_data_q[294]
  PIN i_data_q[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.1850 0.0000 890.2350 0.2200 ;
    END
  END i_data_q[293]
  PIN i_data_q[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.9850 0.0000 890.0350 0.2200 ;
    END
  END i_data_q[292]
  PIN i_data_q[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.7850 0.0000 889.8350 0.2200 ;
    END
  END i_data_q[291]
  PIN i_data_q[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.5850 0.0000 889.6350 0.2200 ;
    END
  END i_data_q[290]
  PIN i_data_q[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.1850 0.0000 889.2350 0.2200 ;
    END
  END i_data_q[289]
  PIN i_data_q[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.9850 0.0000 889.0350 0.2200 ;
    END
  END i_data_q[288]
  PIN i_data_q[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.7850 0.0000 888.8350 0.2200 ;
    END
  END i_data_q[287]
  PIN i_data_q[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.5850 0.0000 888.6350 0.2200 ;
    END
  END i_data_q[286]
  PIN i_data_q[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.3850 0.0000 888.4350 0.2200 ;
    END
  END i_data_q[285]
  PIN i_data_q[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.1850 0.0000 888.2350 0.2200 ;
    END
  END i_data_q[284]
  PIN i_data_q[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.9850 0.0000 888.0350 0.2200 ;
    END
  END i_data_q[283]
  PIN i_data_q[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.7850 0.0000 887.8350 0.2200 ;
    END
  END i_data_q[282]
  PIN i_data_q[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.5850 0.0000 887.6350 0.2200 ;
    END
  END i_data_q[281]
  PIN i_data_q[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.3850 0.0000 887.4350 0.2200 ;
    END
  END i_data_q[280]
  PIN i_data_q[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.9850 0.0000 887.0350 0.2200 ;
    END
  END i_data_q[279]
  PIN i_data_q[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.7850 0.0000 886.8350 0.2200 ;
    END
  END i_data_q[278]
  PIN i_data_q[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.5850 0.0000 886.6350 0.2200 ;
    END
  END i_data_q[277]
  PIN i_data_q[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.3850 0.0000 886.4350 0.2200 ;
    END
  END i_data_q[276]
  PIN i_data_q[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.1850 0.0000 886.2350 0.2200 ;
    END
  END i_data_q[275]
  PIN i_data_q[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.9850 0.0000 886.0350 0.2200 ;
    END
  END i_data_q[274]
  PIN i_data_q[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.7850 0.0000 885.8350 0.2200 ;
    END
  END i_data_q[273]
  PIN i_data_q[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.5850 0.0000 885.6350 0.2200 ;
    END
  END i_data_q[272]
  PIN i_data_q[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.3850 0.0000 885.4350 0.2200 ;
    END
  END i_data_q[271]
  PIN i_data_q[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.1850 0.0000 885.2350 0.2200 ;
    END
  END i_data_q[270]
  PIN i_data_q[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.7850 0.0000 884.8350 0.2200 ;
    END
  END i_data_q[269]
  PIN i_data_q[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.5850 0.0000 884.6350 0.2200 ;
    END
  END i_data_q[268]
  PIN i_data_q[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.3850 0.0000 884.4350 0.2200 ;
    END
  END i_data_q[267]
  PIN i_data_q[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.1850 0.0000 884.2350 0.2200 ;
    END
  END i_data_q[266]
  PIN i_data_q[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.9850 0.0000 884.0350 0.2200 ;
    END
  END i_data_q[265]
  PIN i_data_q[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.7850 0.0000 883.8350 0.2200 ;
    END
  END i_data_q[264]
  PIN i_data_q[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.5850 0.0000 883.6350 0.2200 ;
    END
  END i_data_q[263]
  PIN i_data_q[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.3850 0.0000 883.4350 0.2200 ;
    END
  END i_data_q[262]
  PIN i_data_q[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.1850 0.0000 883.2350 0.2200 ;
    END
  END i_data_q[261]
  PIN i_data_q[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.9850 0.0000 883.0350 0.2200 ;
    END
  END i_data_q[260]
  PIN i_data_q[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.5850 0.0000 882.6350 0.2200 ;
    END
  END i_data_q[259]
  PIN i_data_q[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.3850 0.0000 882.4350 0.2200 ;
    END
  END i_data_q[258]
  PIN i_data_q[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.1850 0.0000 882.2350 0.2200 ;
    END
  END i_data_q[257]
  PIN i_data_q[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.9850 0.0000 882.0350 0.2200 ;
    END
  END i_data_q[256]
  PIN i_data_q[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.7850 0.0000 881.8350 0.2200 ;
    END
  END i_data_q[255]
  PIN i_data_q[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.5850 0.0000 881.6350 0.2200 ;
    END
  END i_data_q[254]
  PIN i_data_q[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.3850 0.0000 881.4350 0.2200 ;
    END
  END i_data_q[253]
  PIN i_data_q[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.1850 0.0000 881.2350 0.2200 ;
    END
  END i_data_q[252]
  PIN i_data_q[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.9850 0.0000 881.0350 0.2200 ;
    END
  END i_data_q[251]
  PIN i_data_q[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.7850 0.0000 880.8350 0.2200 ;
    END
  END i_data_q[250]
  PIN i_data_q[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.3850 0.0000 880.4350 0.2200 ;
    END
  END i_data_q[249]
  PIN i_data_q[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.1850 0.0000 880.2350 0.2200 ;
    END
  END i_data_q[248]
  PIN i_data_q[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.9850 0.0000 880.0350 0.2200 ;
    END
  END i_data_q[247]
  PIN i_data_q[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.7850 0.0000 879.8350 0.2200 ;
    END
  END i_data_q[246]
  PIN i_data_q[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.5850 0.0000 879.6350 0.2200 ;
    END
  END i_data_q[245]
  PIN i_data_q[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.3850 0.0000 879.4350 0.2200 ;
    END
  END i_data_q[244]
  PIN i_data_q[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.1850 0.0000 879.2350 0.2200 ;
    END
  END i_data_q[243]
  PIN i_data_q[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.9850 0.0000 879.0350 0.2200 ;
    END
  END i_data_q[242]
  PIN i_data_q[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.7850 0.0000 878.8350 0.2200 ;
    END
  END i_data_q[241]
  PIN i_data_q[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.5850 0.0000 878.6350 0.2200 ;
    END
  END i_data_q[240]
  PIN i_data_q[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.1850 0.0000 878.2350 0.2200 ;
    END
  END i_data_q[239]
  PIN i_data_q[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 877.9850 0.0000 878.0350 0.2200 ;
    END
  END i_data_q[238]
  PIN i_data_q[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 877.7850 0.0000 877.8350 0.2200 ;
    END
  END i_data_q[237]
  PIN i_data_q[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 874.0850 0.0000 874.1350 0.2200 ;
    END
  END i_data_q[236]
  PIN i_data_q[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.8850 0.0000 873.9350 0.2200 ;
    END
  END i_data_q[235]
  PIN i_data_q[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.6850 0.0000 873.7350 0.2200 ;
    END
  END i_data_q[234]
  PIN i_data_q[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.4850 0.0000 873.5350 0.2200 ;
    END
  END i_data_q[233]
  PIN i_data_q[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.2850 0.0000 873.3350 0.2200 ;
    END
  END i_data_q[232]
  PIN i_data_q[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.0850 0.0000 873.1350 0.2200 ;
    END
  END i_data_q[231]
  PIN i_data_q[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.8850 0.0000 872.9350 0.2200 ;
    END
  END i_data_q[230]
  PIN i_data_q[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.4850 0.0000 872.5350 0.2200 ;
    END
  END i_data_q[229]
  PIN i_data_q[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.2850 0.0000 872.3350 0.2200 ;
    END
  END i_data_q[228]
  PIN i_data_q[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.0850 0.0000 872.1350 0.2200 ;
    END
  END i_data_q[227]
  PIN i_data_q[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.8850 0.0000 871.9350 0.2200 ;
    END
  END i_data_q[226]
  PIN i_data_q[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.6850 0.0000 871.7350 0.2200 ;
    END
  END i_data_q[225]
  PIN i_data_q[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.4850 0.0000 871.5350 0.2200 ;
    END
  END i_data_q[224]
  PIN i_data_q[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.2850 0.0000 871.3350 0.2200 ;
    END
  END i_data_q[223]
  PIN i_data_q[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.0850 0.0000 871.1350 0.2200 ;
    END
  END i_data_q[222]
  PIN i_data_q[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.8850 0.0000 870.9350 0.2200 ;
    END
  END i_data_q[221]
  PIN i_data_q[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.6850 0.0000 870.7350 0.2200 ;
    END
  END i_data_q[220]
  PIN i_data_q[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.2850 0.0000 870.3350 0.2200 ;
    END
  END i_data_q[219]
  PIN i_data_q[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.0850 0.0000 870.1350 0.2200 ;
    END
  END i_data_q[218]
  PIN i_data_q[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.8850 0.0000 869.9350 0.2200 ;
    END
  END i_data_q[217]
  PIN i_data_q[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.6850 0.0000 869.7350 0.2200 ;
    END
  END i_data_q[216]
  PIN i_data_q[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.4850 0.0000 869.5350 0.2200 ;
    END
  END i_data_q[215]
  PIN i_data_q[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.2850 0.0000 869.3350 0.2200 ;
    END
  END i_data_q[214]
  PIN i_data_q[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.0850 0.0000 869.1350 0.2200 ;
    END
  END i_data_q[213]
  PIN i_data_q[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.8850 0.0000 868.9350 0.2200 ;
    END
  END i_data_q[212]
  PIN i_data_q[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.6850 0.0000 868.7350 0.2200 ;
    END
  END i_data_q[211]
  PIN i_data_q[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.4850 0.0000 868.5350 0.2200 ;
    END
  END i_data_q[210]
  PIN i_data_q[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.0850 0.0000 868.1350 0.2200 ;
    END
  END i_data_q[209]
  PIN i_data_q[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.8850 0.0000 867.9350 0.2200 ;
    END
  END i_data_q[208]
  PIN i_data_q[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.6850 0.0000 867.7350 0.2200 ;
    END
  END i_data_q[207]
  PIN i_data_q[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.4850 0.0000 867.5350 0.2200 ;
    END
  END i_data_q[206]
  PIN i_data_q[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.2850 0.0000 867.3350 0.2200 ;
    END
  END i_data_q[205]
  PIN i_data_q[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.0850 0.0000 867.1350 0.2200 ;
    END
  END i_data_q[204]
  PIN i_data_q[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.8850 0.0000 866.9350 0.2200 ;
    END
  END i_data_q[203]
  PIN i_data_q[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.6850 0.0000 866.7350 0.2200 ;
    END
  END i_data_q[202]
  PIN i_data_q[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.4850 0.0000 866.5350 0.2200 ;
    END
  END i_data_q[201]
  PIN i_data_q[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.2850 0.0000 866.3350 0.2200 ;
    END
  END i_data_q[200]
  PIN i_data_q[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.6850 0.0000 865.7350 0.2200 ;
    END
  END i_data_q[199]
  PIN i_data_q[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.4850 0.0000 865.5350 0.2200 ;
    END
  END i_data_q[198]
  PIN i_data_q[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.2850 0.0000 865.3350 0.2200 ;
    END
  END i_data_q[197]
  PIN i_data_q[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.0850 0.0000 865.1350 0.2200 ;
    END
  END i_data_q[196]
  PIN i_data_q[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.8850 0.0000 864.9350 0.2200 ;
    END
  END i_data_q[195]
  PIN i_data_q[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.6850 0.0000 864.7350 0.2200 ;
    END
  END i_data_q[194]
  PIN i_data_q[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.4850 0.0000 864.5350 0.2200 ;
    END
  END i_data_q[193]
  PIN i_data_q[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.2850 0.0000 864.3350 0.2200 ;
    END
  END i_data_q[192]
  PIN i_data_q[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.0850 0.0000 864.1350 0.2200 ;
    END
  END i_data_q[191]
  PIN i_data_q[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.8850 0.0000 863.9350 0.2200 ;
    END
  END i_data_q[190]
  PIN i_data_q[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.4850 0.0000 863.5350 0.2200 ;
    END
  END i_data_q[189]
  PIN i_data_q[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.2850 0.0000 863.3350 0.2200 ;
    END
  END i_data_q[188]
  PIN i_data_q[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.0850 0.0000 863.1350 0.2200 ;
    END
  END i_data_q[187]
  PIN i_data_q[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.8850 0.0000 862.9350 0.2200 ;
    END
  END i_data_q[186]
  PIN i_data_q[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.6850 0.0000 862.7350 0.2200 ;
    END
  END i_data_q[185]
  PIN i_data_q[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.4850 0.0000 862.5350 0.2200 ;
    END
  END i_data_q[184]
  PIN i_data_q[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.2850 0.0000 862.3350 0.2200 ;
    END
  END i_data_q[183]
  PIN i_data_q[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.0850 0.0000 862.1350 0.2200 ;
    END
  END i_data_q[182]
  PIN i_data_q[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.8850 0.0000 861.9350 0.2200 ;
    END
  END i_data_q[181]
  PIN i_data_q[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.6850 0.0000 861.7350 0.2200 ;
    END
  END i_data_q[180]
  PIN i_data_q[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.2850 0.0000 861.3350 0.2200 ;
    END
  END i_data_q[179]
  PIN i_data_q[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.0850 0.0000 861.1350 0.2200 ;
    END
  END i_data_q[178]
  PIN i_data_q[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.8850 0.0000 860.9350 0.2200 ;
    END
  END i_data_q[177]
  PIN i_data_q[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.6850 0.0000 860.7350 0.2200 ;
    END
  END i_data_q[176]
  PIN i_data_q[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.4850 0.0000 860.5350 0.2200 ;
    END
  END i_data_q[175]
  PIN i_data_q[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.2850 0.0000 860.3350 0.2200 ;
    END
  END i_data_q[174]
  PIN i_data_q[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.0850 0.0000 860.1350 0.2200 ;
    END
  END i_data_q[173]
  PIN i_data_q[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.8850 0.0000 859.9350 0.2200 ;
    END
  END i_data_q[172]
  PIN i_data_q[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.6850 0.0000 859.7350 0.2200 ;
    END
  END i_data_q[171]
  PIN i_data_q[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.4850 0.0000 859.5350 0.2200 ;
    END
  END i_data_q[170]
  PIN i_data_q[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.0850 0.0000 859.1350 0.2200 ;
    END
  END i_data_q[169]
  PIN i_data_q[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.8850 0.0000 858.9350 0.2200 ;
    END
  END i_data_q[168]
  PIN i_data_q[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.6850 0.0000 858.7350 0.2200 ;
    END
  END i_data_q[167]
  PIN i_data_q[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.4850 0.0000 858.5350 0.2200 ;
    END
  END i_data_q[166]
  PIN i_data_q[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.2850 0.0000 858.3350 0.2200 ;
    END
  END i_data_q[165]
  PIN i_data_q[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.0850 0.0000 858.1350 0.2200 ;
    END
  END i_data_q[164]
  PIN i_data_q[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.8850 0.0000 857.9350 0.2200 ;
    END
  END i_data_q[163]
  PIN i_data_q[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.6850 0.0000 857.7350 0.2200 ;
    END
  END i_data_q[162]
  PIN i_data_q[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.4850 0.0000 857.5350 0.2200 ;
    END
  END i_data_q[161]
  PIN i_data_q[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.2850 0.0000 857.3350 0.2200 ;
    END
  END i_data_q[160]
  PIN i_data_q[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.8850 0.0000 856.9350 0.2200 ;
    END
  END i_data_q[159]
  PIN i_data_q[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.6850 0.0000 856.7350 0.2200 ;
    END
  END i_data_q[158]
  PIN i_data_q[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.4850 0.0000 856.5350 0.2200 ;
    END
  END i_data_q[157]
  PIN i_data_q[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.2850 0.0000 856.3350 0.2200 ;
    END
  END i_data_q[156]
  PIN i_data_q[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.0850 0.0000 856.1350 0.2200 ;
    END
  END i_data_q[155]
  PIN i_data_q[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.8850 0.0000 855.9350 0.2200 ;
    END
  END i_data_q[154]
  PIN i_data_q[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.6850 0.0000 855.7350 0.2200 ;
    END
  END i_data_q[153]
  PIN i_data_q[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.4850 0.0000 855.5350 0.2200 ;
    END
  END i_data_q[152]
  PIN i_data_q[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.2850 0.0000 855.3350 0.2200 ;
    END
  END i_data_q[151]
  PIN i_data_q[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.0850 0.0000 855.1350 0.2200 ;
    END
  END i_data_q[150]
  PIN i_data_q[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.6850 0.0000 854.7350 0.2200 ;
    END
  END i_data_q[149]
  PIN i_data_q[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.4850 0.0000 854.5350 0.2200 ;
    END
  END i_data_q[148]
  PIN i_data_q[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.2850 0.0000 854.3350 0.2200 ;
    END
  END i_data_q[147]
  PIN i_data_q[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.0850 0.0000 854.1350 0.2200 ;
    END
  END i_data_q[146]
  PIN i_data_q[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.8850 0.0000 853.9350 0.2200 ;
    END
  END i_data_q[145]
  PIN i_data_q[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.6850 0.0000 853.7350 0.2200 ;
    END
  END i_data_q[144]
  PIN i_data_q[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.4850 0.0000 853.5350 0.2200 ;
    END
  END i_data_q[143]
  PIN i_data_q[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.7850 0.0000 849.8350 0.2200 ;
    END
  END i_data_q[142]
  PIN i_data_q[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.5850 0.0000 849.6350 0.2200 ;
    END
  END i_data_q[141]
  PIN i_data_q[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.3850 0.0000 849.4350 0.2200 ;
    END
  END i_data_q[140]
  PIN i_data_q[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.9850 0.0000 849.0350 0.2200 ;
    END
  END i_data_q[139]
  PIN i_data_q[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.7850 0.0000 848.8350 0.2200 ;
    END
  END i_data_q[138]
  PIN i_data_q[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.5850 0.0000 848.6350 0.2200 ;
    END
  END i_data_q[137]
  PIN i_data_q[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.3850 0.0000 848.4350 0.2200 ;
    END
  END i_data_q[136]
  PIN i_data_q[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.1850 0.0000 848.2350 0.2200 ;
    END
  END i_data_q[135]
  PIN i_data_q[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.9850 0.0000 848.0350 0.2200 ;
    END
  END i_data_q[134]
  PIN i_data_q[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.7850 0.0000 847.8350 0.2200 ;
    END
  END i_data_q[133]
  PIN i_data_q[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.5850 0.0000 847.6350 0.2200 ;
    END
  END i_data_q[132]
  PIN i_data_q[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.3850 0.0000 847.4350 0.2200 ;
    END
  END i_data_q[131]
  PIN i_data_q[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.1850 0.0000 847.2350 0.2200 ;
    END
  END i_data_q[130]
  PIN i_data_q[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.7850 0.0000 846.8350 0.2200 ;
    END
  END i_data_q[129]
  PIN i_data_q[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.5850 0.0000 846.6350 0.2200 ;
    END
  END i_data_q[128]
  PIN i_data_q[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.3850 0.0000 846.4350 0.2200 ;
    END
  END i_data_q[127]
  PIN i_data_q[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.1850 0.0000 846.2350 0.2200 ;
    END
  END i_data_q[126]
  PIN i_data_q[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.9850 0.0000 846.0350 0.2200 ;
    END
  END i_data_q[125]
  PIN i_data_q[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.7850 0.0000 845.8350 0.2200 ;
    END
  END i_data_q[124]
  PIN i_data_q[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.5850 0.0000 845.6350 0.2200 ;
    END
  END i_data_q[123]
  PIN i_data_q[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.3850 0.0000 845.4350 0.2200 ;
    END
  END i_data_q[122]
  PIN i_data_q[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.1850 0.0000 845.2350 0.2200 ;
    END
  END i_data_q[121]
  PIN i_data_q[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.9850 0.0000 845.0350 0.2200 ;
    END
  END i_data_q[120]
  PIN i_data_q[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.5850 0.0000 844.6350 0.2200 ;
    END
  END i_data_q[119]
  PIN i_data_q[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.3850 0.0000 844.4350 0.2200 ;
    END
  END i_data_q[118]
  PIN i_data_q[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.1850 0.0000 844.2350 0.2200 ;
    END
  END i_data_q[117]
  PIN i_data_q[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.9850 0.0000 844.0350 0.2200 ;
    END
  END i_data_q[116]
  PIN i_data_q[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.7850 0.0000 843.8350 0.2200 ;
    END
  END i_data_q[115]
  PIN i_data_q[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.5850 0.0000 843.6350 0.2200 ;
    END
  END i_data_q[114]
  PIN i_data_q[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.3850 0.0000 843.4350 0.2200 ;
    END
  END i_data_q[113]
  PIN i_data_q[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.1850 0.0000 843.2350 0.2200 ;
    END
  END i_data_q[112]
  PIN i_data_q[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.9850 0.0000 843.0350 0.2200 ;
    END
  END i_data_q[111]
  PIN i_data_q[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.7850 0.0000 842.8350 0.2200 ;
    END
  END i_data_q[110]
  PIN i_data_q[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.3850 0.0000 842.4350 0.2200 ;
    END
  END i_data_q[109]
  PIN i_data_q[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.1850 0.0000 842.2350 0.2200 ;
    END
  END i_data_q[108]
  PIN i_data_q[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.9850 0.0000 842.0350 0.2200 ;
    END
  END i_data_q[107]
  PIN i_data_q[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.7850 0.0000 841.8350 0.2200 ;
    END
  END i_data_q[106]
  PIN i_data_q[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.5850 0.0000 841.6350 0.2200 ;
    END
  END i_data_q[105]
  PIN i_data_q[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.3850 0.0000 841.4350 0.2200 ;
    END
  END i_data_q[104]
  PIN i_data_q[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.1850 0.0000 841.2350 0.2200 ;
    END
  END i_data_q[103]
  PIN i_data_q[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.9850 0.0000 841.0350 0.2200 ;
    END
  END i_data_q[102]
  PIN i_data_q[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.7850 0.0000 840.8350 0.2200 ;
    END
  END i_data_q[101]
  PIN i_data_q[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.5850 0.0000 840.6350 0.2200 ;
    END
  END i_data_q[100]
  PIN i_data_q[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.5850 0.0000 976.6350 0.2200 ;
    END
  END i_data_q[99]
  PIN i_data_q[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.3850 0.0000 976.4350 0.2200 ;
    END
  END i_data_q[98]
  PIN i_data_q[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.1850 0.0000 976.2350 0.2200 ;
    END
  END i_data_q[97]
  PIN i_data_q[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.9850 0.0000 976.0350 0.2200 ;
    END
  END i_data_q[96]
  PIN i_data_q[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.7850 0.0000 975.8350 0.2200 ;
    END
  END i_data_q[95]
  PIN i_data_q[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.5850 0.0000 975.6350 0.2200 ;
    END
  END i_data_q[94]
  PIN i_data_q[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.3850 0.0000 975.4350 0.2200 ;
    END
  END i_data_q[93]
  PIN i_data_q[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.1850 0.0000 975.2350 0.2200 ;
    END
  END i_data_q[92]
  PIN i_data_q[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.9850 0.0000 975.0350 0.2200 ;
    END
  END i_data_q[91]
  PIN i_data_q[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.7850 0.0000 974.8350 0.2200 ;
    END
  END i_data_q[90]
  PIN i_data_q[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.3850 0.0000 974.4350 0.2200 ;
    END
  END i_data_q[89]
  PIN i_data_q[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.1850 0.0000 974.2350 0.2200 ;
    END
  END i_data_q[88]
  PIN i_data_q[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 970.3850 0.0000 970.4350 0.2200 ;
    END
  END i_data_q[87]
  PIN i_data_q[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 970.1850 0.0000 970.2350 0.2200 ;
    END
  END i_data_q[86]
  PIN i_data_q[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.9850 0.0000 970.0350 0.2200 ;
    END
  END i_data_q[85]
  PIN i_data_q[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.7850 0.0000 969.8350 0.2200 ;
    END
  END i_data_q[84]
  PIN i_data_q[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.5850 0.0000 969.6350 0.2200 ;
    END
  END i_data_q[83]
  PIN i_data_q[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.3850 0.0000 969.4350 0.2200 ;
    END
  END i_data_q[82]
  PIN i_data_q[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.1850 0.0000 969.2350 0.2200 ;
    END
  END i_data_q[81]
  PIN i_data_q[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.9850 0.0000 969.0350 0.2200 ;
    END
  END i_data_q[80]
  PIN i_data_q[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.5850 0.0000 968.6350 0.2200 ;
    END
  END i_data_q[79]
  PIN i_data_q[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.3850 0.0000 968.4350 0.2200 ;
    END
  END i_data_q[78]
  PIN i_data_q[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.1850 0.0000 968.2350 0.2200 ;
    END
  END i_data_q[77]
  PIN i_data_q[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.9850 0.0000 968.0350 0.2200 ;
    END
  END i_data_q[76]
  PIN i_data_q[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.7850 0.0000 967.8350 0.2200 ;
    END
  END i_data_q[75]
  PIN i_data_q[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.5850 0.0000 967.6350 0.2200 ;
    END
  END i_data_q[74]
  PIN i_data_q[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.3850 0.0000 967.4350 0.2200 ;
    END
  END i_data_q[73]
  PIN i_data_q[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.1850 0.0000 967.2350 0.2200 ;
    END
  END i_data_q[72]
  PIN i_data_q[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.9850 0.0000 967.0350 0.2200 ;
    END
  END i_data_q[71]
  PIN i_data_q[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.7850 0.0000 966.8350 0.2200 ;
    END
  END i_data_q[70]
  PIN i_data_q[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.3850 0.0000 966.4350 0.2200 ;
    END
  END i_data_q[69]
  PIN i_data_q[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.1850 0.0000 966.2350 0.2200 ;
    END
  END i_data_q[68]
  PIN i_data_q[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.9850 0.0000 966.0350 0.2200 ;
    END
  END i_data_q[67]
  PIN i_data_q[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.7850 0.0000 965.8350 0.2200 ;
    END
  END i_data_q[66]
  PIN i_data_q[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.5850 0.0000 965.6350 0.2200 ;
    END
  END i_data_q[65]
  PIN i_data_q[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.3850 0.0000 965.4350 0.2200 ;
    END
  END i_data_q[64]
  PIN i_data_q[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.1850 0.0000 965.2350 0.2200 ;
    END
  END i_data_q[63]
  PIN i_data_q[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.9850 0.0000 965.0350 0.2200 ;
    END
  END i_data_q[62]
  PIN i_data_q[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.7850 0.0000 964.8350 0.2200 ;
    END
  END i_data_q[61]
  PIN i_data_q[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.5850 0.0000 964.6350 0.2200 ;
    END
  END i_data_q[60]
  PIN i_data_q[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.1850 0.0000 964.2350 0.2200 ;
    END
  END i_data_q[59]
  PIN i_data_q[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.9850 0.0000 964.0350 0.2200 ;
    END
  END i_data_q[58]
  PIN i_data_q[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.7850 0.0000 963.8350 0.2200 ;
    END
  END i_data_q[57]
  PIN i_data_q[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.3850 0.0000 962.4350 0.2200 ;
    END
  END i_data_q[56]
  PIN i_data_q[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.1850 0.0000 960.2350 0.2200 ;
    END
  END i_data_q[55]
  PIN i_data_q[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.9850 0.0000 958.0350 0.2200 ;
    END
  END i_data_q[54]
  PIN i_data_q[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.7850 0.0000 955.8350 0.2200 ;
    END
  END i_data_q[53]
  PIN i_data_q[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.5850 0.0000 953.6350 0.2200 ;
    END
  END i_data_q[52]
  PIN i_data_q[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.3850 0.0000 951.4350 0.2200 ;
    END
  END i_data_q[51]
  PIN i_data_q[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.5850 0.0000 945.6350 0.2200 ;
    END
  END i_data_q[50]
  PIN i_data_q[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.1850 0.0000 943.2350 0.2200 ;
    END
  END i_data_q[49]
  PIN i_data_q[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.9850 0.0000 941.0350 0.2200 ;
    END
  END i_data_q[48]
  PIN i_data_q[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.7850 0.0000 938.8350 0.2200 ;
    END
  END i_data_q[47]
  PIN i_data_q[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.5850 0.0000 936.6350 0.2200 ;
    END
  END i_data_q[46]
  PIN i_data_q[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.3850 0.0000 934.4350 0.2200 ;
    END
  END i_data_q[45]
  PIN i_data_q[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.1850 0.0000 932.2350 0.2200 ;
    END
  END i_data_q[44]
  PIN i_data_q[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.9850 0.0000 930.0350 0.2200 ;
    END
  END i_data_q[43]
  PIN i_data_q[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.7850 0.0000 927.8350 0.2200 ;
    END
  END i_data_q[42]
  PIN i_data_q[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.9850 0.0000 922.0350 0.2200 ;
    END
  END i_data_q[41]
  PIN i_data_q[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.7850 0.0000 919.8350 0.2200 ;
    END
  END i_data_q[40]
  PIN i_data_q[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.3850 0.0000 917.4350 0.2200 ;
    END
  END i_data_q[39]
  PIN i_data_q[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.1850 0.0000 915.2350 0.2200 ;
    END
  END i_data_q[38]
  PIN i_data_q[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.9850 0.0000 913.0350 0.2200 ;
    END
  END i_data_q[37]
  PIN i_data_q[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.7850 0.0000 910.8350 0.2200 ;
    END
  END i_data_q[36]
  PIN i_data_q[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.5850 0.0000 908.6350 0.2200 ;
    END
  END i_data_q[35]
  PIN i_data_q[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.3850 0.0000 906.4350 0.2200 ;
    END
  END i_data_q[34]
  PIN i_data_q[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.1850 0.0000 904.2350 0.2200 ;
    END
  END i_data_q[33]
  PIN i_data_q[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 898.3850 0.0000 898.4350 0.2200 ;
    END
  END i_data_q[32]
  PIN i_data_q[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.1850 0.0000 896.2350 0.2200 ;
    END
  END i_data_q[31]
  PIN i_data_q[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.9850 0.0000 894.0350 0.2200 ;
    END
  END i_data_q[30]
  PIN i_data_q[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.5850 0.0000 891.6350 0.2200 ;
    END
  END i_data_q[29]
  PIN i_data_q[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.3850 0.0000 889.4350 0.2200 ;
    END
  END i_data_q[28]
  PIN i_data_q[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.1850 0.0000 887.2350 0.2200 ;
    END
  END i_data_q[27]
  PIN i_data_q[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.9850 0.0000 885.0350 0.2200 ;
    END
  END i_data_q[26]
  PIN i_data_q[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.7850 0.0000 882.8350 0.2200 ;
    END
  END i_data_q[25]
  PIN i_data_q[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.5850 0.0000 880.6350 0.2200 ;
    END
  END i_data_q[24]
  PIN i_data_q[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.3850 0.0000 878.4350 0.2200 ;
    END
  END i_data_q[23]
  PIN i_data_q[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.6850 0.0000 872.7350 0.2200 ;
    END
  END i_data_q[22]
  PIN i_data_q[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.4850 0.0000 870.5350 0.2200 ;
    END
  END i_data_q[21]
  PIN i_data_q[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.2850 0.0000 868.3350 0.2200 ;
    END
  END i_data_q[20]
  PIN i_data_q[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.8850 0.0000 865.9350 0.2200 ;
    END
  END i_data_q[19]
  PIN i_data_q[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.6850 0.0000 863.7350 0.2200 ;
    END
  END i_data_q[18]
  PIN i_data_q[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.4850 0.0000 861.5350 0.2200 ;
    END
  END i_data_q[17]
  PIN i_data_q[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.2850 0.0000 859.3350 0.2200 ;
    END
  END i_data_q[16]
  PIN i_data_q[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.0850 0.0000 857.1350 0.2200 ;
    END
  END i_data_q[15]
  PIN i_data_q[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.8850 0.0000 854.9350 0.2200 ;
    END
  END i_data_q[14]
  PIN i_data_q[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.1850 0.0000 849.2350 0.2200 ;
    END
  END i_data_q[13]
  PIN i_data_q[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.9850 0.0000 847.0350 0.2200 ;
    END
  END i_data_q[12]
  PIN i_data_q[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.7850 0.0000 844.8350 0.2200 ;
    END
  END i_data_q[11]
  PIN i_data_q[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.5850 0.0000 842.6350 0.2200 ;
    END
  END i_data_q[10]
  PIN i_data_q[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.7850 0.0000 976.8350 0.2200 ;
    END
  END i_data_q[9]
  PIN i_data_q[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.5850 0.0000 974.6350 0.2200 ;
    END
  END i_data_q[8]
  PIN i_data_q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.7850 0.0000 968.8350 0.2200 ;
    END
  END i_data_q[7]
  PIN i_data_q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.5850 0.0000 966.6350 0.2200 ;
    END
  END i_data_q[6]
  PIN i_data_q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.3850 0.0000 964.4350 0.2200 ;
    END
  END i_data_q[5]
  PIN i_data_q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.3850 0.0000 943.4350 0.2200 ;
    END
  END i_data_q[4]
  PIN i_data_q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.5850 0.0000 917.6350 0.2200 ;
    END
  END i_data_q[3]
  PIN i_data_q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.7850 0.0000 891.8350 0.2200 ;
    END
  END i_data_q[2]
  PIN i_data_q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.0850 0.0000 866.1350 0.2200 ;
    END
  END i_data_q[1]
  PIN i_data_q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.3850 0.0000 840.4350 0.2200 ;
    END
  END i_data_q[0]
  PIN o_fo_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.2850 640.5800 1701.3350 640.8000 ;
    END
  END o_fo_valid
  PIN o_fo_value[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.6850 640.5800 1703.7350 640.8000 ;
    END
  END o_fo_value[14]
  PIN o_fo_value[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 159.8250 1704.3000 159.8750 ;
    END
  END o_fo_value[13]
  PIN o_fo_value[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 191.0250 1704.3000 191.0750 ;
    END
  END o_fo_value[12]
  PIN o_fo_value[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 207.8250 1704.3000 207.8750 ;
    END
  END o_fo_value[11]
  PIN o_fo_value[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 160.5250 1704.3000 160.5750 ;
    END
  END o_fo_value[10]
  PIN o_fo_value[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 163.4250 1704.3000 163.4750 ;
    END
  END o_fo_value[9]
  PIN o_fo_value[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.6850 640.5800 1703.7350 640.8000 ;
    END
  END o_fo_value[8]
  PIN o_fo_value[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.4850 640.5800 1703.5350 640.8000 ;
    END
  END o_fo_value[7]
  PIN o_fo_value[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.4850 640.5800 1703.5350 640.8000 ;
    END
  END o_fo_value[6]
  PIN o_fo_value[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.2850 640.5800 1703.3350 640.8000 ;
    END
  END o_fo_value[5]
  PIN o_fo_value[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.2850 640.5800 1703.3350 640.8000 ;
    END
  END o_fo_value[4]
  PIN o_fo_value[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1703.2100 640.4000 1703.3100 640.8000 ;
    END
  END o_fo_value[3]
  PIN o_fo_value[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.0850 640.5800 1703.1350 640.8000 ;
    END
  END o_fo_value[2]
  PIN o_fo_value[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.0850 640.5800 1703.1350 640.8000 ;
    END
  END o_fo_value[1]
  PIN o_fo_value[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.8850 640.5800 1702.9350 640.8000 ;
    END
  END o_fo_value[0]
  PIN sc_cpren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 3.3250 0.2200 3.3750 ;
    END
  END sc_cpren
  PIN sc_spren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 1.4250 0.2200 1.4750 ;
    END
  END sc_spren
  PIN sc_sen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4850 0.0000 0.5350 0.2200 ;
    END
  END sc_sen
  PIN sc_di0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 51.6850 0.0000 51.7350 0.2200 ;
    END
  END sc_di0
  PIN sc_do0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3850 0.0000 1.4350 0.2200 ;
    END
  END sc_do0
  PIN sc_di1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.6850 0.0000 51.7350 0.2200 ;
    END
  END sc_di1
  PIN sc_do1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.2850 0.0000 2.3350 0.2200 ;
    END
  END sc_do1
  PIN sc_di2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 115.1250 0.2200 115.1750 ;
    END
  END sc_di2
  PIN sc_do2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7850 0.0000 0.8350 0.2200 ;
    END
  END sc_do2
  PIN sc_di3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 272.6250 0.2200 272.6750 ;
    END
  END sc_di3
  PIN sc_do3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.6850 0.0000 2.7350 0.2200 ;
    END
  END sc_do3
  PIN sc_di4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 430.1250 0.2200 430.1750 ;
    END
  END sc_di4
  PIN sc_do4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8.4850 0.0000 8.5350 0.2200 ;
    END
  END sc_do4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER IA ;
        RECT 1427.9020 0.0000 1434.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1451.9020 0.0000 1458.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1331.9020 0.0000 1338.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1355.9020 0.0000 1362.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1379.9020 0.0000 1386.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1403.9020 0.0000 1410.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 920.7980 0.0000 927.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 944.7980 0.0000 951.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 968.7980 0.0000 975.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 992.7980 0.0000 999.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1016.7980 0.0000 1023.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1040.7980 0.0000 1047.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 629.6940 0.0000 636.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 509.6940 0.0000 516.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 533.6940 0.0000 540.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 557.6940 0.0000 564.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 581.6940 0.0000 588.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 605.6940 0.0000 612.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 146.5900 0.0000 153.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 170.5900 0.0000 177.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 194.5900 0.0000 201.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 218.5900 0.0000 225.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 98.5900 0.0000 105.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 122.5900 0.0000 129.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1597.4520 640.4000 1604.4520 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1597.4520 0.0000 1604.4520 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1621.7620 640.4000 1628.7620 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1621.7620 0.0000 1628.7620 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1646.0720 640.4000 1653.0720 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1646.0720 0.0000 1653.0720 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1573.1420 640.4000 1580.1420 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1573.1420 0.0000 1580.1420 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1500.2120 640.4000 1507.2120 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1500.2120 0.0000 1507.2120 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1524.5220 640.4000 1531.5220 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1524.5220 0.0000 1531.5220 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1548.8320 640.4000 1555.8320 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1548.8320 0.0000 1555.8320 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1475.9020 640.4000 1482.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1475.9020 0.0000 1482.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1307.9020 640.4000 1314.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1307.9020 0.0000 1314.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1259.2780 640.4000 1266.2780 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1259.2780 0.0000 1266.2780 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1283.5880 640.4000 1290.5880 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1283.5880 0.0000 1290.5880 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1186.3480 640.4000 1193.3480 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1186.3480 0.0000 1193.3480 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1210.6580 640.4000 1217.6580 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1210.6580 0.0000 1217.6580 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1234.9680 640.4000 1241.9680 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1234.9680 0.0000 1241.9680 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1113.4180 640.4000 1120.4180 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1113.4180 0.0000 1120.4180 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1137.7280 640.4000 1144.7280 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1137.7280 0.0000 1144.7280 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1162.0380 640.4000 1169.0380 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1162.0380 0.0000 1169.0380 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1064.7980 640.4000 1071.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1064.7980 0.0000 1071.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1089.1080 640.4000 1096.1080 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1089.1080 0.0000 1096.1080 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 896.7980 640.4000 903.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 896.7980 0.0000 903.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 872.4840 640.4000 879.4840 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 872.4840 0.0000 879.4840 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 848.1740 640.4000 855.1740 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 848.1740 0.0000 855.1740 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 775.2440 640.4000 782.2440 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 775.2440 0.0000 782.2440 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 799.5540 640.4000 806.5540 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 799.5540 0.0000 806.5540 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 823.8640 640.4000 830.8640 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 823.8640 0.0000 830.8640 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 702.3140 640.4000 709.3140 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 702.3140 0.0000 709.3140 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 726.6240 640.4000 733.6240 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 726.6240 0.0000 733.6240 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 750.9340 640.4000 757.9340 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 750.9340 0.0000 757.9340 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 653.6940 640.4000 660.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 653.6940 0.0000 660.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 678.0040 640.4000 685.0040 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 678.0040 0.0000 685.0040 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 485.6940 640.4000 492.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 485.6940 0.0000 492.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 461.3800 640.4000 468.3800 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 461.3800 0.0000 468.3800 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 388.4500 640.4000 395.4500 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 388.4500 0.0000 395.4500 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 412.7600 640.4000 419.7600 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 412.7600 0.0000 419.7600 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 437.0700 640.4000 444.0700 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 437.0700 0.0000 444.0700 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 291.2100 640.4000 298.2100 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 291.2100 0.0000 298.2100 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 315.5200 640.4000 322.5200 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 315.5200 0.0000 322.5200 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 339.8300 640.4000 346.8300 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 339.8300 0.0000 346.8300 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 364.1400 640.4000 371.1400 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 364.1400 0.0000 371.1400 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 242.5900 640.4000 249.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 242.5900 0.0000 249.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 266.9000 640.4000 273.9000 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 266.9000 0.0000 273.9000 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 74.5900 640.4000 81.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 74.5900 0.0000 81.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 50.2760 640.4000 57.2760 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 50.2760 0.0000 57.2760 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 25.9660 640.4000 32.9660 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 25.9660 0.0000 32.9660 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1.6560 640.4000 8.6560 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1.6560 0.0000 8.6560 0.4000 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 640.7330 0.0500 640.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 640.7330 1704.3000 640.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 638.3330 0.0500 638.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 638.3330 1704.3000 638.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 633.5330 0.0500 633.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 633.5330 1704.3000 633.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 635.9330 0.0500 636.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 635.9330 1704.3000 636.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 628.7330 0.0500 628.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 628.7330 1704.3000 628.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 631.1330 0.0500 631.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 631.1330 1704.3000 631.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 623.9330 0.0500 624.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 623.9330 1704.3000 624.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 626.3330 0.0500 626.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 626.3330 1704.3000 626.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 621.5330 0.0500 621.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 621.5330 1704.3000 621.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 618.0960 0.4000 625.0960 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 618.0960 1704.3000 625.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 616.7330 0.0500 616.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 616.7330 1704.3000 616.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 619.1330 0.0500 619.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 619.1330 1704.3000 619.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 611.9330 0.0500 612.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 611.9330 1704.3000 612.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 614.3330 0.0500 614.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 614.3330 1704.3000 614.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 607.1330 0.0500 607.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 607.1330 1704.3000 607.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 609.5330 0.0500 609.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 609.5330 1704.3000 609.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 604.7330 0.0500 604.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 604.7330 1704.3000 604.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 602.3330 0.0500 602.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 602.3330 1704.3000 602.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 597.5330 0.0500 597.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 597.5330 1704.3000 597.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 599.9330 0.0500 600.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 599.9330 1704.3000 600.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 594.4680 0.4000 601.4680 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 594.4680 1704.3000 601.4680 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 592.7330 0.0500 592.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 592.7330 1704.3000 592.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 595.1330 0.0500 595.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 595.1330 1704.3000 595.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 587.9330 0.0500 588.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 587.9330 1704.3000 588.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 590.3330 0.0500 590.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 590.3330 1704.3000 590.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 583.1330 0.0500 583.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 583.1330 1704.3000 583.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 585.5330 0.0500 585.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 585.5330 1704.3000 585.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 578.3330 0.0500 578.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 578.3330 1704.3000 578.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 580.7330 0.0500 580.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 580.7330 1704.3000 580.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 570.8400 0.4000 577.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 570.8400 1704.3000 577.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 573.5330 0.0500 573.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 573.5330 1704.3000 573.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 575.9330 0.0500 576.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 575.9330 1704.3000 576.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 571.1330 0.0500 571.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 571.1330 1704.3000 571.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 566.3330 0.0500 566.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 566.3330 1704.3000 566.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 568.7330 0.0500 568.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 568.7330 1704.3000 568.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 561.5330 0.0500 561.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 561.5330 1704.3000 561.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 563.9330 0.0500 564.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 563.9330 1704.3000 564.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 556.7330 0.0500 556.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 556.7330 1704.3000 556.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 559.1330 0.0500 559.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 559.1330 1704.3000 559.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 506.3330 0.0500 506.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 506.3330 1704.3000 506.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 498.8400 0.4000 505.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 498.8400 1704.3000 505.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 503.9330 0.0500 504.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 503.9330 1704.3000 504.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 501.5330 0.0500 501.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 501.5330 1704.3000 501.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 499.1330 0.0500 499.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 499.1330 1704.3000 499.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 496.7330 0.0500 496.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 496.7330 1704.3000 496.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 494.3330 0.0500 494.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 494.3330 1704.3000 494.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 491.9330 0.0500 492.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 491.9330 1704.3000 492.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 489.5330 0.0500 489.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 489.5330 1704.3000 489.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 487.1330 0.0500 487.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 487.1330 1704.3000 487.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 484.7330 0.0500 484.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 484.7330 1704.3000 484.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 482.3330 0.0500 482.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 482.3330 1704.3000 482.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 479.9330 0.0500 480.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 479.9330 1704.3000 480.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 477.5330 0.0500 477.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 477.5330 1704.3000 477.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 475.2040 0.4000 482.2040 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 475.2040 1704.3000 482.2040 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 475.1330 0.0500 475.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 475.1330 1704.3000 475.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 472.7330 0.0500 472.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 472.7330 1704.3000 472.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 465.5330 0.0500 465.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 465.5330 1704.3000 465.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 467.9330 0.0500 468.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 467.9330 1704.3000 468.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 470.3330 0.0500 470.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 470.3330 1704.3000 470.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 460.7330 0.0500 460.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 460.7330 1704.3000 460.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 463.1330 0.0500 463.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 463.1330 1704.3000 463.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 455.9330 0.0500 456.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 455.9330 1704.3000 456.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 458.3330 0.0500 458.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 458.3330 1704.3000 458.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 451.5760 0.4000 458.5760 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 451.5760 1704.3000 458.5760 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 451.1330 0.0500 451.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 451.1330 1704.3000 451.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 453.5330 0.0500 453.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 453.5330 1704.3000 453.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 446.3330 0.0500 446.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 446.3330 1704.3000 446.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 448.7330 0.0500 448.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 448.7330 1704.3000 448.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 441.5330 0.0500 441.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 441.5330 1704.3000 441.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 443.9330 0.0500 444.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 443.9330 1704.3000 444.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 436.7330 0.0500 436.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 436.7330 1704.3000 436.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 439.1330 0.0500 439.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 439.1330 1704.3000 439.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 431.9330 0.0500 432.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 431.9330 1704.3000 432.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 434.3330 0.0500 434.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 434.3330 1704.3000 434.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 427.9480 0.4000 434.9480 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 427.9480 1704.3000 434.9480 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 427.1330 0.0500 427.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 427.1330 1704.3000 427.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 429.5330 0.0500 429.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 429.5330 1704.3000 429.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 422.3330 0.0500 422.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 422.3330 1704.3000 422.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 424.7330 0.0500 424.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 424.7330 1704.3000 424.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 417.5330 0.0500 417.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 417.5330 1704.3000 417.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 419.9330 0.0500 420.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 419.9330 1704.3000 420.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 415.1330 0.0500 415.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 415.1330 1704.3000 415.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 410.3330 0.0500 410.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 410.3330 1704.3000 410.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 412.7330 0.0500 412.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 412.7330 1704.3000 412.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 405.5330 0.0500 405.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 405.5330 1704.3000 405.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 407.9330 0.0500 408.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 407.9330 1704.3000 408.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 404.3200 0.4000 411.3200 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 404.3200 1704.3000 411.3200 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 400.7330 0.0500 400.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 400.7330 1704.3000 400.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 403.1330 0.0500 403.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 403.1330 1704.3000 403.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 395.9330 0.0500 396.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 395.9330 1704.3000 396.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 398.3330 0.0500 398.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 398.3330 1704.3000 398.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 391.1330 0.0500 391.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 391.1330 1704.3000 391.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 393.5330 0.0500 393.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 393.5330 1704.3000 393.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 386.3330 0.0500 386.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 386.3330 1704.3000 386.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 388.7330 0.0500 388.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 388.7330 1704.3000 388.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 380.6920 0.4000 387.6920 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 380.6920 1704.3000 387.6920 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 381.5330 0.0500 381.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 381.5330 1704.3000 381.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 383.9330 0.0500 384.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 383.9330 1704.3000 384.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 376.7330 0.0500 376.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 376.7330 1704.3000 376.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 379.1330 0.0500 379.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 379.1330 1704.3000 379.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 371.9330 0.0500 372.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 371.9330 1704.3000 372.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 374.3330 0.0500 374.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 374.3330 1704.3000 374.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 367.1330 0.0500 367.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 367.1330 1704.3000 367.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 369.5330 0.0500 369.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 369.5330 1704.3000 369.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 364.7330 0.0500 364.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 364.7330 1704.3000 364.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 359.9330 0.0500 360.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 359.9330 1704.3000 360.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 362.3330 0.0500 362.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 362.3330 1704.3000 362.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 357.0640 0.4000 364.0640 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 357.0640 1704.3000 364.0640 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 357.5330 0.0500 357.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 357.5330 1704.3000 357.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 355.1330 0.0500 355.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 355.1330 1704.3000 355.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 350.3330 0.0500 350.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 350.3330 1704.3000 350.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 352.7330 0.0500 352.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 352.7330 1704.3000 352.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 345.5330 0.0500 345.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 345.5330 1704.3000 345.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 347.9330 0.0500 348.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 347.9330 1704.3000 348.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 340.7330 0.0500 340.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 340.7330 1704.3000 340.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 343.1330 0.0500 343.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 343.1330 1704.3000 343.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 338.3330 0.0500 338.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 338.3330 1704.3000 338.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 335.9330 0.0500 336.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 335.9330 1704.3000 336.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 333.4360 0.4000 340.4360 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 333.4360 1704.3000 340.4360 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 331.1330 0.0500 331.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 331.1330 1704.3000 331.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 333.5330 0.0500 333.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 333.5330 1704.3000 333.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 326.3330 0.0500 326.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 326.3330 1704.3000 326.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 328.7330 0.0500 328.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 328.7330 1704.3000 328.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 321.5330 0.0500 321.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 321.5330 1704.3000 321.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 323.9330 0.0500 324.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 323.9330 1704.3000 324.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 316.7330 0.0500 316.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 316.7330 1704.3000 316.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 319.1330 0.0500 319.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 319.1330 1704.3000 319.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 309.8080 0.4000 316.8080 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 309.8080 1704.3000 316.8080 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 309.5330 0.0500 309.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 309.5330 1704.3000 309.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 311.9330 0.0500 312.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 311.9330 1704.3000 312.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 314.3330 0.0500 314.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 314.3330 1704.3000 314.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 304.7330 0.0500 304.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 304.7330 1704.3000 304.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 307.1330 0.0500 307.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 307.1330 1704.3000 307.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 299.9330 0.0500 300.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 299.9330 1704.3000 300.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 302.3330 0.0500 302.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 302.3330 1704.3000 302.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 295.1330 0.0500 295.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 295.1330 1704.3000 295.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 297.5330 0.0500 297.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 297.5330 1704.3000 297.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 290.3330 0.0500 290.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 290.3330 1704.3000 290.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 292.7330 0.0500 292.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 292.7330 1704.3000 292.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 286.1800 0.4000 293.1800 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 286.1800 1704.3000 293.1800 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 285.5330 0.0500 285.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 285.5330 1704.3000 285.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 287.9330 0.0500 288.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 287.9330 1704.3000 288.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 280.7330 0.0500 280.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 280.7330 1704.3000 280.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 283.1330 0.0500 283.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 283.1330 1704.3000 283.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 275.9330 0.0500 276.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 275.9330 1704.3000 276.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 278.3330 0.0500 278.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 278.3330 1704.3000 278.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 271.1330 0.0500 271.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 271.1330 1704.3000 271.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 273.5330 0.0500 273.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 273.5330 1704.3000 273.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 266.3330 0.0500 266.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 266.3330 1704.3000 266.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 268.7330 0.0500 268.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 268.7330 1704.3000 268.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 262.5520 0.4000 269.5520 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 262.5520 1704.3000 269.5520 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 261.5330 0.0500 261.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 261.5330 1704.3000 261.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 263.9330 0.0500 264.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 263.9330 1704.3000 264.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 259.1330 0.0500 259.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 259.1330 1704.3000 259.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 254.3330 0.0500 254.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 254.3330 1704.3000 254.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 256.7330 0.0500 256.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 256.7330 1704.3000 256.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 249.5330 0.0500 249.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 249.5330 1704.3000 249.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 251.9330 0.0500 252.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 251.9330 1704.3000 252.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 244.7330 0.0500 244.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 244.7330 1704.3000 244.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 247.1330 0.0500 247.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 247.1330 1704.3000 247.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 238.9240 0.4000 245.9240 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 238.9240 1704.3000 245.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 239.9330 0.0500 240.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 239.9330 1704.3000 240.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 242.3330 0.0500 242.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 242.3330 1704.3000 242.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 235.1330 0.0500 235.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 235.1330 1704.3000 235.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 237.5330 0.0500 237.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 237.5330 1704.3000 237.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 230.3330 0.0500 230.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 230.3330 1704.3000 230.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 232.7330 0.0500 232.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 232.7330 1704.3000 232.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 225.5330 0.0500 225.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 225.5330 1704.3000 225.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 227.9330 0.0500 228.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 227.9330 1704.3000 228.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 220.7330 0.0500 220.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 220.7330 1704.3000 220.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 223.1330 0.0500 223.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 223.1330 1704.3000 223.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 215.2960 0.4000 222.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 215.2960 1704.3000 222.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 215.9330 0.0500 216.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 215.9330 1704.3000 216.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 218.3330 0.0500 218.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 218.3330 1704.3000 218.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 211.1330 0.0500 211.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 211.1330 1704.3000 211.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 213.5330 0.0500 213.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 213.5330 1704.3000 213.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 208.7330 0.0500 208.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 208.7330 1704.3000 208.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 206.3330 0.0500 206.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 206.3330 1704.3000 206.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 203.9330 0.0500 204.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 203.9330 1704.3000 204.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 201.5330 0.0500 201.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 201.5330 1704.3000 201.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 148.7330 0.0500 148.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 148.7330 1704.3000 148.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 151.1330 0.0500 151.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 151.1330 1704.3000 151.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 146.3330 0.0500 146.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 146.3330 1704.3000 146.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 143.9330 0.0500 144.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 143.9330 1704.3000 144.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 143.2960 0.4000 150.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 143.2960 1704.3000 150.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 139.1330 0.0500 139.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 139.1330 1704.3000 139.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 141.5330 0.0500 141.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 141.5330 1704.3000 141.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 136.7330 0.0500 136.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 136.7330 1704.3000 136.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 134.3330 0.0500 134.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 134.3330 1704.3000 134.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 131.9330 0.0500 132.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 131.9330 1704.3000 132.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 129.5330 0.0500 129.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 129.5330 1704.3000 129.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 127.1330 0.0500 127.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 127.1330 1704.3000 127.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 124.7330 0.0500 124.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 124.7330 1704.3000 124.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 119.6600 0.4000 126.6600 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 119.6600 1704.3000 126.6600 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 122.3330 0.0500 122.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 122.3330 1704.3000 122.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 119.9330 0.0500 120.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 119.9330 1704.3000 120.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 117.5330 0.0500 117.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 117.5330 1704.3000 117.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 115.1330 0.0500 115.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 115.1330 1704.3000 115.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 112.7330 0.0500 112.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 112.7330 1704.3000 112.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 110.3330 0.0500 110.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 110.3330 1704.3000 110.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 107.9330 0.0500 108.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 107.9330 1704.3000 108.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 105.5330 0.0500 105.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 105.5330 1704.3000 105.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 103.1330 0.0500 103.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 103.1330 1704.3000 103.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 100.7330 0.0500 100.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 100.7330 1704.3000 100.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 98.3330 0.0500 98.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 98.3330 1704.3000 98.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 96.0320 0.4000 103.0320 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 96.0320 1704.3000 103.0320 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 95.9330 0.0500 96.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 95.9330 1704.3000 96.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 93.5330 0.0500 93.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 93.5330 1704.3000 93.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 91.1330 0.0500 91.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 91.1330 1704.3000 91.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 88.7330 0.0500 88.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 88.7330 1704.3000 88.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 86.3330 0.0500 86.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 86.3330 1704.3000 86.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 83.9330 0.0500 84.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 83.9330 1704.3000 84.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 81.5330 0.0500 81.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 81.5330 1704.3000 81.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 79.1330 0.0500 79.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 79.1330 1704.3000 79.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.7330 0.0500 76.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 76.7330 1704.3000 76.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 74.3330 0.0500 74.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 74.3330 1704.3000 74.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 72.4040 0.4000 79.4040 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 72.4040 1704.3000 79.4040 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 71.9330 0.0500 72.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 71.9330 1704.3000 72.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 69.5330 0.0500 69.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 69.5330 1704.3000 69.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 67.1330 0.0500 67.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 67.1330 1704.3000 67.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 64.7330 0.0500 64.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 64.7330 1704.3000 64.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 62.3330 0.0500 62.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 62.3330 1704.3000 62.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 59.9330 0.0500 60.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 59.9330 1704.3000 60.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 57.5330 0.0500 57.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 57.5330 1704.3000 57.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 55.1330 0.0500 55.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 55.1330 1704.3000 55.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 52.7330 0.0500 52.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 52.7330 1704.3000 52.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 48.7760 0.4000 55.7760 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 48.7760 1704.3000 55.7760 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 50.3330 0.0500 50.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 50.3330 1704.3000 50.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 47.9330 0.0500 48.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 47.9330 1704.3000 48.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 45.5330 0.0500 45.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 45.5330 1704.3000 45.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 43.1330 0.0500 43.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 43.1330 1704.3000 43.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 40.7330 0.0500 40.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 40.7330 1704.3000 40.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 38.3330 0.0500 38.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 38.3330 1704.3000 38.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 35.9330 0.0500 36.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 35.9330 1704.3000 36.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 33.5330 0.0500 33.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 33.5330 1704.3000 33.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 31.1330 0.0500 31.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 31.1330 1704.3000 31.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.7330 0.0500 28.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 28.7330 1704.3000 28.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 25.1480 0.4000 32.1480 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 25.1480 1704.3000 32.1480 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 26.3330 0.0500 26.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 26.3330 1704.3000 26.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 23.9330 0.0500 24.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 23.9330 1704.3000 24.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 21.5330 0.0500 21.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 21.5330 1704.3000 21.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 19.1330 0.0500 19.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 19.1330 1704.3000 19.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7330 0.0500 16.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 16.7330 1704.3000 16.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 14.3330 0.0500 14.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 14.3330 1704.3000 14.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 11.9330 0.0500 12.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 11.9330 1704.3000 12.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.5330 0.0500 9.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 9.5330 1704.3000 9.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 7.1330 0.0500 7.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 7.1330 1704.3000 7.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 4.7330 0.0500 4.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 4.7330 1704.3000 4.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 2.3330 0.0500 2.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 2.3330 1704.3000 2.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 1.5200 0.4000 8.5200 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 1.5200 1704.3000 8.5200 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 -0.0670 0.0500 0.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 -0.0670 1704.3000 0.0670 ;
    END
    PORT
      LAYER IA ;
        RECT 1694.6920 640.4000 1701.6920 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1694.6920 0.0000 1701.6920 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1670.3820 640.4000 1677.3820 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1670.3820 0.0000 1677.3820 0.4000 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 191.2960 0.4000 198.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 167.2960 0.4000 174.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 153.5330 0.0500 153.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 155.9330 0.0500 156.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 158.3330 0.0500 158.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 160.7330 0.0500 160.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 163.1330 0.0500 163.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 165.5330 0.0500 165.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 167.9330 0.0500 168.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 170.3330 0.0500 170.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 172.7330 0.0500 172.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 175.1330 0.0500 175.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 177.5330 0.0500 177.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 179.9330 0.0500 180.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 182.3330 0.0500 182.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 184.7330 0.0500 184.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 187.1330 0.0500 187.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 189.5330 0.0500 189.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 191.9330 0.0500 192.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 194.3330 0.0500 194.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 196.7330 0.0500 196.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 199.1330 0.0500 199.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 546.8400 0.4000 553.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 522.8400 0.4000 529.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 508.7330 0.0500 508.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 511.1330 0.0500 511.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 513.5330 0.0500 513.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 515.9330 0.0500 516.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 518.3330 0.0500 518.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 520.7330 0.0500 520.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 523.1330 0.0500 523.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 525.5330 0.0500 525.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 527.9330 0.0500 528.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 530.3330 0.0500 530.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 532.7330 0.0500 532.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 535.1330 0.0500 535.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 537.5330 0.0500 537.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 539.9330 0.0500 540.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 542.3330 0.0500 542.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 544.7330 0.0500 544.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 547.1330 0.0500 547.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 549.5330 0.0500 549.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 551.9330 0.0500 552.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 554.3330 0.0500 554.4670 ;
    END
    PORT
      LAYER IA ;
        RECT 122.5900 640.4000 129.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 98.5900 640.4000 105.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 218.5900 640.4000 225.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 194.5900 640.4000 201.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 170.5900 640.4000 177.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 146.5900 640.4000 153.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 605.6940 640.4000 612.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 581.6940 640.4000 588.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 557.6940 640.4000 564.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 533.6940 640.4000 540.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 509.6940 640.4000 516.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 629.6940 640.4000 636.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 920.7980 640.4000 927.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1040.7980 640.4000 1047.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1016.7980 640.4000 1023.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 992.7980 640.4000 999.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 968.7980 640.4000 975.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 944.7980 640.4000 951.7980 640.8000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 153.5330 1704.3000 153.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 155.9330 1704.3000 156.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 158.3330 1704.3000 158.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 160.7330 1704.3000 160.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 163.1330 1704.3000 163.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 167.2960 1704.3000 174.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 165.5330 1704.3000 165.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 167.9330 1704.3000 168.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 170.3330 1704.3000 170.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 172.7330 1704.3000 172.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 175.1330 1704.3000 175.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 177.5330 1704.3000 177.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 179.9330 1704.3000 180.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 182.3330 1704.3000 182.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 191.2960 1704.3000 198.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 184.7330 1704.3000 184.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 187.1330 1704.3000 187.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 189.5330 1704.3000 189.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 191.9330 1704.3000 192.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 194.3330 1704.3000 194.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 196.7330 1704.3000 196.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 199.1330 1704.3000 199.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 508.7330 1704.3000 508.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 511.1330 1704.3000 511.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 513.5330 1704.3000 513.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 515.9330 1704.3000 516.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 518.3330 1704.3000 518.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 520.7330 1704.3000 520.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 523.1330 1704.3000 523.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 525.5330 1704.3000 525.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 522.8400 1704.3000 529.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 546.8400 1704.3000 553.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 527.9330 1704.3000 528.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 530.3330 1704.3000 530.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 532.7330 1704.3000 532.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 535.1330 1704.3000 535.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 537.5330 1704.3000 537.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 539.9330 1704.3000 540.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 542.3330 1704.3000 542.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 544.7330 1704.3000 544.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 547.1330 1704.3000 547.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 549.5330 1704.3000 549.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 551.9330 1704.3000 552.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 554.3330 1704.3000 554.4670 ;
    END
    PORT
      LAYER IA ;
        RECT 1403.9020 640.4000 1410.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1379.9020 640.4000 1386.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1355.9020 640.4000 1362.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1331.9020 640.4000 1338.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1451.9020 640.4000 1458.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1427.9020 640.4000 1434.9020 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1700.3000 491.8400 1704.3000 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1700.3000 136.2960 1704.3000 166.2960 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER IA ;
        RECT 1439.9020 0.0000 1446.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1415.9020 0.0000 1422.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1319.9020 0.0000 1326.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1343.9020 0.0000 1350.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1367.9020 0.0000 1374.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1391.9020 0.0000 1398.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 908.7980 0.0000 915.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 932.7980 0.0000 939.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 956.7980 0.0000 963.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 980.7980 0.0000 987.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1004.7980 0.0000 1011.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1028.7980 0.0000 1035.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 617.6940 0.0000 624.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 497.6940 0.0000 504.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 521.6940 0.0000 528.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 545.6940 0.0000 552.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 569.6940 0.0000 576.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 593.6940 0.0000 600.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 134.5900 0.0000 141.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 158.5900 0.0000 165.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 182.5900 0.0000 189.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 206.5900 0.0000 213.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 86.5900 0.0000 93.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 110.5900 0.0000 117.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1585.2970 640.4000 1592.2970 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1585.2970 0.0000 1592.2970 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1609.6070 640.4000 1616.6070 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1609.6070 0.0000 1616.6070 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1633.9170 640.4000 1640.9170 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1633.9170 0.0000 1640.9170 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1512.3670 640.4000 1519.3670 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1512.3670 0.0000 1519.3670 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1536.6770 640.4000 1543.6770 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1536.6770 0.0000 1543.6770 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1560.9870 640.4000 1567.9870 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1560.9870 0.0000 1567.9870 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1463.9020 640.4000 1470.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1463.9020 0.0000 1470.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1488.0570 640.4000 1495.0570 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1488.0570 0.0000 1495.0570 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1271.4330 640.4000 1278.4330 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1271.4330 0.0000 1278.4330 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1295.7430 640.4000 1302.7430 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1295.7430 0.0000 1302.7430 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1198.5030 640.4000 1205.5030 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1198.5030 0.0000 1205.5030 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1222.8130 640.4000 1229.8130 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1222.8130 0.0000 1229.8130 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1247.1230 640.4000 1254.1230 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1247.1230 0.0000 1254.1230 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1174.1930 640.4000 1181.1930 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1174.1930 0.0000 1181.1930 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1101.2630 640.4000 1108.2630 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1101.2630 0.0000 1108.2630 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1125.5730 640.4000 1132.5730 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1125.5730 0.0000 1132.5730 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1149.8830 640.4000 1156.8830 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1149.8830 0.0000 1156.8830 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1052.7980 640.4000 1059.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1052.7980 0.0000 1059.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1076.9530 640.4000 1083.9530 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1076.9530 0.0000 1083.9530 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 860.3290 640.4000 867.3290 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 860.3290 0.0000 867.3290 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 884.6390 640.4000 891.6390 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 884.6390 0.0000 891.6390 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 787.3990 640.4000 794.3990 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 787.3990 0.0000 794.3990 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 811.7090 640.4000 818.7090 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 811.7090 0.0000 818.7090 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 836.0190 640.4000 843.0190 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 836.0190 0.0000 843.0190 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 714.4690 640.4000 721.4690 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 714.4690 0.0000 721.4690 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 738.7790 640.4000 745.7790 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 738.7790 0.0000 745.7790 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 763.0890 640.4000 770.0890 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 763.0890 0.0000 770.0890 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 690.1590 640.4000 697.1590 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 690.1590 0.0000 697.1590 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 641.6940 640.4000 648.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 641.6940 0.0000 648.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 665.8490 640.4000 672.8490 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 665.8490 0.0000 672.8490 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 473.5350 640.4000 480.5350 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 473.5350 0.0000 480.5350 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 449.2250 640.4000 456.2250 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 449.2250 0.0000 456.2250 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 376.2950 640.4000 383.2950 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 376.2950 0.0000 383.2950 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 400.6050 640.4000 407.6050 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 400.6050 0.0000 407.6050 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 424.9150 640.4000 431.9150 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 424.9150 0.0000 431.9150 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 303.3650 640.4000 310.3650 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 303.3650 0.0000 310.3650 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 327.6750 640.4000 334.6750 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 327.6750 0.0000 334.6750 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 351.9850 640.4000 358.9850 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 351.9850 0.0000 358.9850 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 230.5900 640.4000 237.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 230.5900 0.0000 237.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 254.7450 640.4000 261.7450 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 254.7450 0.0000 261.7450 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 279.0550 640.4000 286.0550 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 279.0550 0.0000 286.0550 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 62.4310 640.4000 69.4310 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 62.4310 0.0000 69.4310 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 13.8110 640.4000 20.8110 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 13.8110 0.0000 20.8110 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 38.1210 640.4000 45.1210 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 38.1210 0.0000 45.1210 0.4000 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 639.5330 0.0500 639.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 639.5330 1704.3000 639.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 637.1330 0.0500 637.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 637.1330 1704.3000 637.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 629.9100 0.4000 636.9100 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 629.9100 1704.3000 636.9100 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 632.3330 0.0500 632.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 632.3330 1704.3000 632.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 634.7330 0.0500 634.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 634.7330 1704.3000 634.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 627.5330 0.0500 627.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 627.5330 1704.3000 627.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 629.9330 0.0500 630.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 629.9330 1704.3000 630.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 622.7330 0.0500 622.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 622.7330 1704.3000 622.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 625.1330 0.0500 625.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 625.1330 1704.3000 625.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 620.3330 0.0500 620.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 620.3330 1704.3000 620.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 617.9330 0.0500 618.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 617.9330 1704.3000 618.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 613.1330 0.0500 613.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 613.1330 1704.3000 613.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 615.5330 0.0500 615.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 615.5330 1704.3000 615.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 608.3330 0.0500 608.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 608.3330 1704.3000 608.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 610.7330 0.0500 610.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 610.7330 1704.3000 610.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 606.2820 0.4000 613.2820 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 606.2820 1704.3000 613.2820 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 603.5330 0.0500 603.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 603.5330 1704.3000 603.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 605.9330 0.0500 606.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 605.9330 1704.3000 606.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 598.7330 0.0500 598.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 598.7330 1704.3000 598.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 601.1330 0.0500 601.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 601.1330 1704.3000 601.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 596.3330 0.0500 596.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 596.3330 1704.3000 596.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 591.5330 0.0500 591.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 591.5330 1704.3000 591.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 593.9330 0.0500 594.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 593.9330 1704.3000 594.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 586.7330 0.0500 586.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 586.7330 1704.3000 586.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 589.1330 0.0500 589.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 589.1330 1704.3000 589.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 582.6540 0.4000 589.6540 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 582.6540 1704.3000 589.6540 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 581.9330 0.0500 582.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 581.9330 1704.3000 582.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 584.3330 0.0500 584.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 584.3330 1704.3000 584.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 577.1330 0.0500 577.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 577.1330 1704.3000 577.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 579.5330 0.0500 579.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 579.5330 1704.3000 579.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 572.3330 0.0500 572.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 572.3330 1704.3000 572.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 574.7330 0.0500 574.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 574.7330 1704.3000 574.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 567.5330 0.0500 567.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 567.5330 1704.3000 567.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 569.9330 0.0500 570.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 569.9330 1704.3000 570.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 562.7330 0.0500 562.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 562.7330 1704.3000 562.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 565.1330 0.0500 565.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 565.1330 1704.3000 565.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 558.8400 0.4000 565.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 558.8400 1704.3000 565.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 557.9330 0.0500 558.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 557.9330 1704.3000 558.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 560.3330 0.0500 560.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 560.3330 1704.3000 560.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 555.5330 0.0500 555.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 555.5330 1704.3000 555.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 505.1330 0.0500 505.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 505.1330 1704.3000 505.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 502.7330 0.0500 502.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 502.7330 1704.3000 502.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 500.3330 0.0500 500.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 500.3330 1704.3000 500.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 497.9330 0.0500 498.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 497.9330 1704.3000 498.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 495.5330 0.0500 495.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 495.5330 1704.3000 495.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 493.1330 0.0500 493.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 493.1330 1704.3000 493.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 490.7330 0.0500 490.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 490.7330 1704.3000 490.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 487.0180 0.4000 494.0180 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 487.0180 1704.3000 494.0180 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 488.3330 0.0500 488.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 488.3330 1704.3000 488.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 485.9330 0.0500 486.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 485.9330 1704.3000 486.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 483.5330 0.0500 483.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 483.5330 1704.3000 483.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 481.1330 0.0500 481.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 481.1330 1704.3000 481.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 478.7330 0.0500 478.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 478.7330 1704.3000 478.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 476.3330 0.0500 476.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 476.3330 1704.3000 476.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 473.9330 0.0500 474.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 473.9330 1704.3000 474.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 471.5330 0.0500 471.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 471.5330 1704.3000 471.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 466.7330 0.0500 466.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 466.7330 1704.3000 466.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 469.1330 0.0500 469.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 469.1330 1704.3000 469.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 463.3900 0.4000 470.3900 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 463.3900 1704.3000 470.3900 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 464.3330 0.0500 464.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 464.3330 1704.3000 464.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 461.9330 0.0500 462.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 461.9330 1704.3000 462.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 459.5330 0.0500 459.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 459.5330 1704.3000 459.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 457.1330 0.0500 457.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 457.1330 1704.3000 457.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 454.7330 0.0500 454.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 454.7330 1704.3000 454.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 452.3330 0.0500 452.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 452.3330 1704.3000 452.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 449.9330 0.0500 450.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 449.9330 1704.3000 450.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 447.5330 0.0500 447.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 447.5330 1704.3000 447.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 439.7620 0.4000 446.7620 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 439.7620 1704.3000 446.7620 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 445.1330 0.0500 445.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 445.1330 1704.3000 445.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 442.7330 0.0500 442.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 442.7330 1704.3000 442.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 440.3330 0.0500 440.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 440.3330 1704.3000 440.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 437.9330 0.0500 438.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 437.9330 1704.3000 438.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 435.5330 0.0500 435.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 435.5330 1704.3000 435.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 433.1330 0.0500 433.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 433.1330 1704.3000 433.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 430.7330 0.0500 430.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 430.7330 1704.3000 430.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 428.3330 0.0500 428.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 428.3330 1704.3000 428.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 425.9330 0.0500 426.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 425.9330 1704.3000 426.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 423.5330 0.0500 423.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 423.5330 1704.3000 423.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 421.1330 0.0500 421.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 421.1330 1704.3000 421.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 416.1340 0.4000 423.1340 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 416.1340 1704.3000 423.1340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 418.7330 0.0500 418.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 418.7330 1704.3000 418.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 416.3330 0.0500 416.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 416.3330 1704.3000 416.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 411.5330 0.0500 411.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 411.5330 1704.3000 411.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 413.9330 0.0500 414.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 413.9330 1704.3000 414.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 409.1330 0.0500 409.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 409.1330 1704.3000 409.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 406.7330 0.0500 406.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 406.7330 1704.3000 406.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 404.3330 0.0500 404.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 404.3330 1704.3000 404.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 401.9330 0.0500 402.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 401.9330 1704.3000 402.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 399.5330 0.0500 399.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 399.5330 1704.3000 399.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 397.1330 0.0500 397.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 397.1330 1704.3000 397.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 392.5060 0.4000 399.5060 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 392.5060 1704.3000 399.5060 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 392.3330 0.0500 392.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 392.3330 1704.3000 392.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 394.7330 0.0500 394.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 394.7330 1704.3000 394.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 389.9330 0.0500 390.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 389.9330 1704.3000 390.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 385.1330 0.0500 385.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 385.1330 1704.3000 385.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 387.5330 0.0500 387.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 387.5330 1704.3000 387.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 380.3330 0.0500 380.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 380.3330 1704.3000 380.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 382.7330 0.0500 382.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 382.7330 1704.3000 382.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 377.9330 0.0500 378.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 377.9330 1704.3000 378.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 375.5330 0.0500 375.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 375.5330 1704.3000 375.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 368.8780 0.4000 375.8780 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 368.8780 1704.3000 375.8780 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 370.7330 0.0500 370.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 370.7330 1704.3000 370.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 373.1330 0.0500 373.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 373.1330 1704.3000 373.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 365.9330 0.0500 366.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 365.9330 1704.3000 366.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 368.3330 0.0500 368.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 368.3330 1704.3000 368.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 361.1330 0.0500 361.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 361.1330 1704.3000 361.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 363.5330 0.0500 363.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 363.5330 1704.3000 363.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 358.7330 0.0500 358.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 358.7330 1704.3000 358.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 356.3330 0.0500 356.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 356.3330 1704.3000 356.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 351.5330 0.0500 351.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 351.5330 1704.3000 351.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 353.9330 0.0500 354.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 353.9330 1704.3000 354.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 345.2500 0.4000 352.2500 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 345.2500 1704.3000 352.2500 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 346.7330 0.0500 346.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 346.7330 1704.3000 346.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 349.1330 0.0500 349.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 349.1330 1704.3000 349.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 341.9330 0.0500 342.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 341.9330 1704.3000 342.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 344.3330 0.0500 344.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 344.3330 1704.3000 344.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 339.5330 0.0500 339.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 339.5330 1704.3000 339.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 334.7330 0.0500 334.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 334.7330 1704.3000 334.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 337.1330 0.0500 337.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 337.1330 1704.3000 337.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 329.9330 0.0500 330.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 329.9330 1704.3000 330.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 332.3330 0.0500 332.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 332.3330 1704.3000 332.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 325.1330 0.0500 325.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 325.1330 1704.3000 325.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 327.5330 0.0500 327.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 327.5330 1704.3000 327.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 321.6220 0.4000 328.6220 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 321.6220 1704.3000 328.6220 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 320.3330 0.0500 320.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 320.3330 1704.3000 320.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 322.7330 0.0500 322.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 322.7330 1704.3000 322.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 315.5330 0.0500 315.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 315.5330 1704.3000 315.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 317.9330 0.0500 318.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 317.9330 1704.3000 318.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 310.7330 0.0500 310.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 310.7330 1704.3000 310.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 313.1330 0.0500 313.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 313.1330 1704.3000 313.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 305.9330 0.0500 306.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 305.9330 1704.3000 306.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 308.3330 0.0500 308.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 308.3330 1704.3000 308.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 297.9940 0.4000 304.9940 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 297.9940 1704.3000 304.9940 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 301.1330 0.0500 301.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 301.1330 1704.3000 301.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 303.5330 0.0500 303.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 303.5330 1704.3000 303.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 296.3330 0.0500 296.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 296.3330 1704.3000 296.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 298.7330 0.0500 298.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 298.7330 1704.3000 298.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 291.5330 0.0500 291.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 291.5330 1704.3000 291.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 293.9330 0.0500 294.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 293.9330 1704.3000 294.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 284.3330 0.0500 284.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 284.3330 1704.3000 284.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 286.7330 0.0500 286.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 286.7330 1704.3000 286.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 289.1330 0.0500 289.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 289.1330 1704.3000 289.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 279.5330 0.0500 279.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 279.5330 1704.3000 279.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 281.9330 0.0500 282.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 281.9330 1704.3000 282.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 274.3660 0.4000 281.3660 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 274.3660 1704.3000 281.3660 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 274.7330 0.0500 274.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 274.7330 1704.3000 274.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 277.1330 0.0500 277.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 277.1330 1704.3000 277.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 269.9330 0.0500 270.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 269.9330 1704.3000 270.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 272.3330 0.0500 272.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 272.3330 1704.3000 272.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 265.1330 0.0500 265.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 265.1330 1704.3000 265.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 267.5330 0.0500 267.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 267.5330 1704.3000 267.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 262.7330 0.0500 262.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 262.7330 1704.3000 262.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 260.3330 0.0500 260.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 260.3330 1704.3000 260.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 255.5330 0.0500 255.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 255.5330 1704.3000 255.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 257.9330 0.0500 258.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 257.9330 1704.3000 258.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 250.7380 0.4000 257.7380 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 250.7380 1704.3000 257.7380 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 250.7330 0.0500 250.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 250.7330 1704.3000 250.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 253.1330 0.0500 253.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 253.1330 1704.3000 253.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 245.9330 0.0500 246.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 245.9330 1704.3000 246.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 248.3330 0.0500 248.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 248.3330 1704.3000 248.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 241.1330 0.0500 241.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 241.1330 1704.3000 241.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 243.5330 0.0500 243.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 243.5330 1704.3000 243.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 236.3330 0.0500 236.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 236.3330 1704.3000 236.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 238.7330 0.0500 238.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 238.7330 1704.3000 238.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 233.9330 0.0500 234.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 233.9330 1704.3000 234.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 227.1100 0.4000 234.1100 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 227.1100 1704.3000 234.1100 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 229.1330 0.0500 229.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 229.1330 1704.3000 229.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 231.5330 0.0500 231.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 231.5330 1704.3000 231.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 224.3330 0.0500 224.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 224.3330 1704.3000 224.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 226.7330 0.0500 226.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 226.7330 1704.3000 226.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 219.5330 0.0500 219.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 219.5330 1704.3000 219.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 221.9330 0.0500 222.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 221.9330 1704.3000 222.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 214.7330 0.0500 214.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 214.7330 1704.3000 214.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 217.1330 0.0500 217.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 217.1330 1704.3000 217.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 209.9330 0.0500 210.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 209.9330 1704.3000 210.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 212.3330 0.0500 212.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 212.3330 1704.3000 212.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 207.5330 0.0500 207.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 207.5330 1704.3000 207.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 205.1330 0.0500 205.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 205.1330 1704.3000 205.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 203.2960 0.4000 210.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 203.2960 1704.3000 210.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 202.7330 0.0500 202.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 202.7330 1704.3000 202.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 200.3330 0.0500 200.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 200.3330 1704.3000 200.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 149.9330 0.0500 150.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 149.9330 1704.3000 150.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 145.1330 0.0500 145.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 145.1330 1704.3000 145.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 147.5330 0.0500 147.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 147.5330 1704.3000 147.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 140.3330 0.0500 140.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 140.3330 1704.3000 140.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 142.7330 0.0500 142.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 142.7330 1704.3000 142.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 137.9330 0.0500 138.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 137.9330 1704.3000 138.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 135.5330 0.0500 135.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 135.5330 1704.3000 135.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 131.4740 0.4000 138.4740 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 131.4740 1704.3000 138.4740 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 133.1330 0.0500 133.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 133.1330 1704.3000 133.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 130.7330 0.0500 130.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 130.7330 1704.3000 130.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 128.3330 0.0500 128.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 128.3330 1704.3000 128.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 125.9330 0.0500 126.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 125.9330 1704.3000 126.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 123.5330 0.0500 123.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 123.5330 1704.3000 123.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 121.1330 0.0500 121.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 121.1330 1704.3000 121.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 118.7330 0.0500 118.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 118.7330 1704.3000 118.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 116.3330 0.0500 116.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 116.3330 1704.3000 116.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 113.9330 0.0500 114.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 113.9330 1704.3000 114.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 107.8460 0.4000 114.8460 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 107.8460 1704.3000 114.8460 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 111.5330 0.0500 111.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 111.5330 1704.3000 111.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 109.1330 0.0500 109.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 109.1330 1704.3000 109.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 106.7330 0.0500 106.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 106.7330 1704.3000 106.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 104.3330 0.0500 104.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 104.3330 1704.3000 104.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 101.9330 0.0500 102.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 101.9330 1704.3000 102.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 99.5330 0.0500 99.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 99.5330 1704.3000 99.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 97.1330 0.0500 97.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 97.1330 1704.3000 97.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 94.7330 0.0500 94.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 94.7330 1704.3000 94.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 92.3330 0.0500 92.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 92.3330 1704.3000 92.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 89.9330 0.0500 90.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 89.9330 1704.3000 90.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 84.2180 0.4000 91.2180 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 84.2180 1704.3000 91.2180 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 87.5330 0.0500 87.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 87.5330 1704.3000 87.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 85.1330 0.0500 85.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 85.1330 1704.3000 85.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 82.7330 0.0500 82.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 82.7330 1704.3000 82.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 80.3330 0.0500 80.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 80.3330 1704.3000 80.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 77.9330 0.0500 78.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 77.9330 1704.3000 78.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 75.5330 0.0500 75.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 75.5330 1704.3000 75.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 73.1330 0.0500 73.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 73.1330 1704.3000 73.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 70.7330 0.0500 70.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 70.7330 1704.3000 70.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 68.3330 0.0500 68.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 68.3330 1704.3000 68.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 65.9330 0.0500 66.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 65.9330 1704.3000 66.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 63.5330 0.0500 63.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 63.5330 1704.3000 63.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 60.5900 0.4000 67.5900 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 60.5900 1704.3000 67.5900 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 61.1330 0.0500 61.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 61.1330 1704.3000 61.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 58.7330 0.0500 58.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 58.7330 1704.3000 58.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 56.3330 0.0500 56.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 56.3330 1704.3000 56.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 53.9330 0.0500 54.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 53.9330 1704.3000 54.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 51.5330 0.0500 51.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 51.5330 1704.3000 51.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 49.1330 0.0500 49.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 49.1330 1704.3000 49.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 46.7330 0.0500 46.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 46.7330 1704.3000 46.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 44.3330 0.0500 44.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 44.3330 1704.3000 44.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 36.9620 0.4000 43.9620 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 36.9620 1704.3000 43.9620 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.9330 0.0500 42.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 41.9330 1704.3000 42.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 39.5330 0.0500 39.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 39.5330 1704.3000 39.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 37.1330 0.0500 37.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 37.1330 1704.3000 37.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 34.7330 0.0500 34.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 34.7330 1704.3000 34.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.3330 0.0500 32.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 32.3330 1704.3000 32.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 29.9330 0.0500 30.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 29.9330 1704.3000 30.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 27.5330 0.0500 27.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 27.5330 1704.3000 27.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.1330 0.0500 25.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 25.1330 1704.3000 25.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 22.7330 0.0500 22.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 22.7330 1704.3000 22.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 20.3330 0.0500 20.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 20.3330 1704.3000 20.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.9330 0.0500 18.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 17.9330 1704.3000 18.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 13.3340 0.4000 20.3340 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 13.3340 1704.3000 20.3340 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 15.5330 0.0500 15.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 15.5330 1704.3000 15.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 13.1330 0.0500 13.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 13.1330 1704.3000 13.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 10.7330 0.0500 10.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 10.7330 1704.3000 10.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 8.3330 0.0500 8.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 8.3330 1704.3000 8.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 5.9330 0.0500 6.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 5.9330 1704.3000 6.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 3.5330 0.0500 3.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 3.5330 1704.3000 3.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 1.1330 0.0500 1.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 1.1330 1704.3000 1.2670 ;
    END
    PORT
      LAYER IA ;
        RECT 1658.2270 640.4000 1665.2270 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1658.2270 0.0000 1665.2270 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1682.5370 640.4000 1689.5370 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1682.5370 0.0000 1689.5370 0.4000 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 179.2960 0.4000 186.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 155.2960 0.4000 162.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 152.3330 0.0500 152.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 154.7330 0.0500 154.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 157.1330 0.0500 157.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 159.5330 0.0500 159.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 161.9330 0.0500 162.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 164.3330 0.0500 164.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 166.7330 0.0500 166.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 169.1330 0.0500 169.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 171.5330 0.0500 171.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 173.9330 0.0500 174.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 176.3330 0.0500 176.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 178.7330 0.0500 178.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 181.1330 0.0500 181.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 183.5330 0.0500 183.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 185.9330 0.0500 186.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 188.3330 0.0500 188.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 190.7330 0.0500 190.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 193.1330 0.0500 193.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 195.5330 0.0500 195.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 197.9330 0.0500 198.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 534.8400 0.4000 541.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 510.8400 0.4000 517.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 507.5330 0.0500 507.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 509.9330 0.0500 510.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 512.3330 0.0500 512.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 514.7330 0.0500 514.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 517.1330 0.0500 517.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 519.5330 0.0500 519.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 521.9330 0.0500 522.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 524.3330 0.0500 524.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 526.7330 0.0500 526.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 529.1330 0.0500 529.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 531.5330 0.0500 531.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 533.9330 0.0500 534.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 536.3330 0.0500 536.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 538.7330 0.0500 538.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 541.1330 0.0500 541.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 543.5330 0.0500 543.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 545.9330 0.0500 546.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 548.3330 0.0500 548.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 550.7330 0.0500 550.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 553.1330 0.0500 553.2670 ;
    END
    PORT
      LAYER IA ;
        RECT 110.5900 640.4000 117.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 86.5900 640.4000 93.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 206.5900 640.4000 213.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 182.5900 640.4000 189.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 158.5900 640.4000 165.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 134.5900 640.4000 141.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 593.6940 640.4000 600.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 569.6940 640.4000 576.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 545.6940 640.4000 552.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 521.6940 640.4000 528.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 497.6940 640.4000 504.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 617.6940 640.4000 624.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 908.7980 640.4000 915.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 932.7980 640.4000 939.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1028.7980 640.4000 1035.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1004.7980 640.4000 1011.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 980.7980 640.4000 987.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 956.7980 640.4000 963.7980 640.8000 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 155.2960 1704.3000 162.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 152.3330 1704.3000 152.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 154.7330 1704.3000 154.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 157.1330 1704.3000 157.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 159.5330 1704.3000 159.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 161.9330 1704.3000 162.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 164.3330 1704.3000 164.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 166.7330 1704.3000 166.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 169.1330 1704.3000 169.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 171.5330 1704.3000 171.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 173.9330 1704.3000 174.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 176.3330 1704.3000 176.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 178.7330 1704.3000 178.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 181.1330 1704.3000 181.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 179.2960 1704.3000 186.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 183.5330 1704.3000 183.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 185.9330 1704.3000 186.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 188.3330 1704.3000 188.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 190.7330 1704.3000 190.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 193.1330 1704.3000 193.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 195.5330 1704.3000 195.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 197.9330 1704.3000 198.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 510.8400 1704.3000 517.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 507.5330 1704.3000 507.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 509.9330 1704.3000 510.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 512.3330 1704.3000 512.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 514.7330 1704.3000 514.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 517.1330 1704.3000 517.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 519.5330 1704.3000 519.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 521.9330 1704.3000 522.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 524.3330 1704.3000 524.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 1703.9000 534.8400 1704.3000 541.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 526.7330 1704.3000 526.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 529.1330 1704.3000 529.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 531.5330 1704.3000 531.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 533.9330 1704.3000 534.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 536.3330 1704.3000 536.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 538.7330 1704.3000 538.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 541.1330 1704.3000 541.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 543.5330 1704.3000 543.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 545.9330 1704.3000 546.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 548.3330 1704.3000 548.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 550.7330 1704.3000 550.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 553.1330 1704.3000 553.2670 ;
    END
    PORT
      LAYER IA ;
        RECT 1391.9020 640.4000 1398.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1367.9020 640.4000 1374.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1343.9020 640.4000 1350.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1319.9020 640.4000 1326.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1415.9020 640.4000 1422.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1439.9020 640.4000 1446.9020 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1700.3000 546.8400 1704.3000 576.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1700.3000 191.2960 1704.3000 221.2960 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 1704.3000 640.8000 ;
    LAYER M2 ;
      RECT 0.2600 640.5230 1704.0400 640.8000 ;
      RECT 0.0000 639.8770 1704.3000 640.5230 ;
      RECT 0.2600 639.3230 1704.0400 639.8770 ;
      RECT 0.0000 638.6770 1704.3000 639.3230 ;
      RECT 0.2600 638.1230 1704.0400 638.6770 ;
      RECT 0.0000 637.4770 1704.3000 638.1230 ;
      RECT 0.2600 636.9230 1704.0400 637.4770 ;
      RECT 0.0000 636.2770 1704.3000 636.9230 ;
      RECT 0.2600 635.7230 1704.0400 636.2770 ;
      RECT 0.0000 635.0770 1704.3000 635.7230 ;
      RECT 0.2600 634.5230 1704.0400 635.0770 ;
      RECT 0.0000 633.8770 1704.3000 634.5230 ;
      RECT 0.2600 633.3230 1704.0400 633.8770 ;
      RECT 0.0000 632.6770 1704.3000 633.3230 ;
      RECT 0.2600 632.1230 1704.0400 632.6770 ;
      RECT 0.0000 631.4770 1704.3000 632.1230 ;
      RECT 0.2600 630.9230 1704.0400 631.4770 ;
      RECT 0.0000 630.2770 1704.3000 630.9230 ;
      RECT 0.2600 629.7230 1704.0400 630.2770 ;
      RECT 0.0000 629.0770 1704.3000 629.7230 ;
      RECT 0.2600 628.5230 1704.0400 629.0770 ;
      RECT 0.0000 627.8770 1704.3000 628.5230 ;
      RECT 0.2600 627.3230 1704.0400 627.8770 ;
      RECT 0.0000 626.6770 1704.3000 627.3230 ;
      RECT 0.2600 626.1230 1704.0400 626.6770 ;
      RECT 0.0000 625.4770 1704.3000 626.1230 ;
      RECT 0.2600 624.9230 1704.0400 625.4770 ;
      RECT 0.0000 624.2770 1704.3000 624.9230 ;
      RECT 0.2600 623.7230 1704.0400 624.2770 ;
      RECT 0.0000 623.0770 1704.3000 623.7230 ;
      RECT 0.2600 622.5230 1704.0400 623.0770 ;
      RECT 0.0000 621.8770 1704.3000 622.5230 ;
      RECT 0.2600 621.3230 1704.0400 621.8770 ;
      RECT 0.0000 620.6770 1704.3000 621.3230 ;
      RECT 0.2600 620.1230 1704.0400 620.6770 ;
      RECT 0.0000 619.4770 1704.3000 620.1230 ;
      RECT 0.2600 618.9230 1704.0400 619.4770 ;
      RECT 0.0000 618.2770 1704.3000 618.9230 ;
      RECT 0.2600 617.7230 1704.0400 618.2770 ;
      RECT 0.0000 617.0770 1704.3000 617.7230 ;
      RECT 0.2600 616.5230 1704.0400 617.0770 ;
      RECT 0.0000 615.8770 1704.3000 616.5230 ;
      RECT 0.2600 615.3230 1704.0400 615.8770 ;
      RECT 0.0000 614.6770 1704.3000 615.3230 ;
      RECT 0.2600 614.1230 1704.0400 614.6770 ;
      RECT 0.0000 613.4770 1704.3000 614.1230 ;
      RECT 0.2600 612.9230 1704.0400 613.4770 ;
      RECT 0.0000 612.2770 1704.3000 612.9230 ;
      RECT 0.2600 611.7230 1704.0400 612.2770 ;
      RECT 0.0000 611.0770 1704.3000 611.7230 ;
      RECT 0.2600 610.5230 1704.0400 611.0770 ;
      RECT 0.0000 609.8770 1704.3000 610.5230 ;
      RECT 0.2600 609.3230 1704.0400 609.8770 ;
      RECT 0.0000 608.6770 1704.3000 609.3230 ;
      RECT 0.2600 608.1230 1704.0400 608.6770 ;
      RECT 0.0000 607.4770 1704.3000 608.1230 ;
      RECT 0.2600 606.9230 1704.0400 607.4770 ;
      RECT 0.0000 606.2770 1704.3000 606.9230 ;
      RECT 0.2600 605.7230 1704.0400 606.2770 ;
      RECT 0.0000 605.0770 1704.3000 605.7230 ;
      RECT 0.2600 604.5230 1704.0400 605.0770 ;
      RECT 0.0000 603.8770 1704.3000 604.5230 ;
      RECT 0.2600 603.3230 1704.0400 603.8770 ;
      RECT 0.0000 602.6770 1704.3000 603.3230 ;
      RECT 0.2600 602.1230 1704.0400 602.6770 ;
      RECT 0.0000 601.4770 1704.3000 602.1230 ;
      RECT 0.2600 600.9230 1704.0400 601.4770 ;
      RECT 0.0000 600.2770 1704.3000 600.9230 ;
      RECT 0.2600 599.7230 1704.0400 600.2770 ;
      RECT 0.0000 599.0770 1704.3000 599.7230 ;
      RECT 0.2600 598.5230 1704.0400 599.0770 ;
      RECT 0.0000 597.8770 1704.3000 598.5230 ;
      RECT 0.2600 597.3230 1704.0400 597.8770 ;
      RECT 0.0000 596.6770 1704.3000 597.3230 ;
      RECT 0.2600 596.1230 1704.0400 596.6770 ;
      RECT 0.0000 595.4770 1704.3000 596.1230 ;
      RECT 0.2600 594.9230 1704.0400 595.4770 ;
      RECT 0.0000 594.2770 1704.3000 594.9230 ;
      RECT 0.2600 593.7230 1704.0400 594.2770 ;
      RECT 0.0000 593.0770 1704.3000 593.7230 ;
      RECT 0.2600 592.5230 1704.0400 593.0770 ;
      RECT 0.0000 591.8770 1704.3000 592.5230 ;
      RECT 0.2600 591.3230 1704.0400 591.8770 ;
      RECT 0.0000 590.6770 1704.3000 591.3230 ;
      RECT 0.2600 590.1230 1704.0400 590.6770 ;
      RECT 0.0000 589.4770 1704.3000 590.1230 ;
      RECT 0.2600 588.9230 1704.0400 589.4770 ;
      RECT 0.0000 588.2770 1704.3000 588.9230 ;
      RECT 0.2600 587.7230 1704.0400 588.2770 ;
      RECT 0.0000 587.0770 1704.3000 587.7230 ;
      RECT 0.2600 586.5230 1704.0400 587.0770 ;
      RECT 0.0000 585.8770 1704.3000 586.5230 ;
      RECT 0.2600 585.3230 1704.0400 585.8770 ;
      RECT 0.0000 584.6770 1704.3000 585.3230 ;
      RECT 0.2600 584.1230 1704.0400 584.6770 ;
      RECT 0.0000 583.4770 1704.3000 584.1230 ;
      RECT 0.2600 582.9230 1704.0400 583.4770 ;
      RECT 0.0000 582.2770 1704.3000 582.9230 ;
      RECT 0.2600 581.7230 1704.0400 582.2770 ;
      RECT 0.0000 581.0770 1704.3000 581.7230 ;
      RECT 0.2600 580.5230 1704.0400 581.0770 ;
      RECT 0.0000 579.8770 1704.3000 580.5230 ;
      RECT 0.2600 579.3230 1704.0400 579.8770 ;
      RECT 0.0000 578.6770 1704.3000 579.3230 ;
      RECT 0.2600 578.1230 1704.0400 578.6770 ;
      RECT 0.0000 577.4770 1704.3000 578.1230 ;
      RECT 0.2600 576.9230 1704.0400 577.4770 ;
      RECT 0.0000 576.2770 1704.3000 576.9230 ;
      RECT 0.2600 575.7230 1704.0400 576.2770 ;
      RECT 0.0000 575.0770 1704.3000 575.7230 ;
      RECT 0.2600 574.5230 1704.0400 575.0770 ;
      RECT 0.0000 573.8770 1704.3000 574.5230 ;
      RECT 0.2600 573.3230 1704.0400 573.8770 ;
      RECT 0.0000 572.6770 1704.3000 573.3230 ;
      RECT 0.2600 572.1230 1704.0400 572.6770 ;
      RECT 0.0000 571.4770 1704.3000 572.1230 ;
      RECT 0.2600 570.9230 1704.0400 571.4770 ;
      RECT 0.0000 570.2770 1704.3000 570.9230 ;
      RECT 0.2600 569.7230 1704.0400 570.2770 ;
      RECT 0.0000 569.0770 1704.3000 569.7230 ;
      RECT 0.2600 568.5230 1704.0400 569.0770 ;
      RECT 0.0000 567.8770 1704.3000 568.5230 ;
      RECT 0.2600 567.3230 1704.0400 567.8770 ;
      RECT 0.0000 566.6770 1704.3000 567.3230 ;
      RECT 0.2600 566.1230 1704.0400 566.6770 ;
      RECT 0.0000 565.4770 1704.3000 566.1230 ;
      RECT 0.2600 564.9230 1704.0400 565.4770 ;
      RECT 0.0000 564.2770 1704.3000 564.9230 ;
      RECT 0.2600 563.7230 1704.0400 564.2770 ;
      RECT 0.0000 563.0770 1704.3000 563.7230 ;
      RECT 0.2600 562.5230 1704.0400 563.0770 ;
      RECT 0.0000 561.8770 1704.3000 562.5230 ;
      RECT 0.2600 561.3230 1704.0400 561.8770 ;
      RECT 0.0000 560.6770 1704.3000 561.3230 ;
      RECT 0.2600 560.1230 1704.0400 560.6770 ;
      RECT 0.0000 559.4770 1704.3000 560.1230 ;
      RECT 0.2600 558.9230 1704.0400 559.4770 ;
      RECT 0.0000 558.2770 1704.3000 558.9230 ;
      RECT 0.2600 557.7230 1704.0400 558.2770 ;
      RECT 0.0000 557.0770 1704.3000 557.7230 ;
      RECT 0.2600 556.5230 1704.0400 557.0770 ;
      RECT 0.0000 555.8770 1704.3000 556.5230 ;
      RECT 0.2600 555.3230 1704.0400 555.8770 ;
      RECT 0.0000 554.6770 1704.3000 555.3230 ;
      RECT 0.2600 554.1230 1704.0400 554.6770 ;
      RECT 0.0000 553.4770 1704.3000 554.1230 ;
      RECT 0.2600 552.9230 1704.0400 553.4770 ;
      RECT 0.0000 552.2770 1704.3000 552.9230 ;
      RECT 0.2600 551.7230 1704.0400 552.2770 ;
      RECT 0.0000 551.0770 1704.3000 551.7230 ;
      RECT 0.2600 550.5230 1704.0400 551.0770 ;
      RECT 0.0000 549.8770 1704.3000 550.5230 ;
      RECT 0.2600 549.3230 1704.0400 549.8770 ;
      RECT 0.0000 548.6770 1704.3000 549.3230 ;
      RECT 0.2600 548.1230 1704.0400 548.6770 ;
      RECT 0.0000 547.4770 1704.3000 548.1230 ;
      RECT 0.2600 546.9230 1704.0400 547.4770 ;
      RECT 0.0000 546.2770 1704.3000 546.9230 ;
      RECT 0.2600 545.7230 1704.0400 546.2770 ;
      RECT 0.0000 545.0770 1704.3000 545.7230 ;
      RECT 0.2600 544.5230 1704.0400 545.0770 ;
      RECT 0.0000 543.8770 1704.3000 544.5230 ;
      RECT 0.2600 543.3230 1704.0400 543.8770 ;
      RECT 0.0000 542.6770 1704.3000 543.3230 ;
      RECT 0.2600 542.1230 1704.0400 542.6770 ;
      RECT 0.0000 541.4770 1704.3000 542.1230 ;
      RECT 0.2600 540.9230 1704.0400 541.4770 ;
      RECT 0.0000 540.2770 1704.3000 540.9230 ;
      RECT 0.2600 539.7230 1704.0400 540.2770 ;
      RECT 0.0000 539.0770 1704.3000 539.7230 ;
      RECT 0.2600 538.5230 1704.0400 539.0770 ;
      RECT 0.0000 537.8770 1704.3000 538.5230 ;
      RECT 0.2600 537.3230 1704.0400 537.8770 ;
      RECT 0.0000 536.6770 1704.3000 537.3230 ;
      RECT 0.2600 536.1230 1704.0400 536.6770 ;
      RECT 0.0000 535.4770 1704.3000 536.1230 ;
      RECT 0.2600 534.9230 1704.0400 535.4770 ;
      RECT 0.0000 534.2770 1704.3000 534.9230 ;
      RECT 0.2600 533.7230 1704.0400 534.2770 ;
      RECT 0.0000 533.0770 1704.3000 533.7230 ;
      RECT 0.2600 532.5230 1704.0400 533.0770 ;
      RECT 0.0000 531.8770 1704.3000 532.5230 ;
      RECT 0.2600 531.3230 1704.0400 531.8770 ;
      RECT 0.0000 530.6770 1704.3000 531.3230 ;
      RECT 0.2600 530.1230 1704.0400 530.6770 ;
      RECT 0.0000 529.4770 1704.3000 530.1230 ;
      RECT 0.2600 528.9230 1704.0400 529.4770 ;
      RECT 0.0000 528.2770 1704.3000 528.9230 ;
      RECT 0.2600 527.7230 1704.0400 528.2770 ;
      RECT 0.0000 527.0770 1704.3000 527.7230 ;
      RECT 0.2600 526.5230 1704.0400 527.0770 ;
      RECT 0.0000 525.8770 1704.3000 526.5230 ;
      RECT 0.2600 525.3230 1704.0400 525.8770 ;
      RECT 0.0000 524.6770 1704.3000 525.3230 ;
      RECT 0.2600 524.1230 1704.0400 524.6770 ;
      RECT 0.0000 523.4770 1704.3000 524.1230 ;
      RECT 0.2600 522.9230 1704.0400 523.4770 ;
      RECT 0.0000 522.2770 1704.3000 522.9230 ;
      RECT 0.2600 521.7230 1704.0400 522.2770 ;
      RECT 0.0000 521.0770 1704.3000 521.7230 ;
      RECT 0.2600 520.5230 1704.0400 521.0770 ;
      RECT 0.0000 519.8770 1704.3000 520.5230 ;
      RECT 0.2600 519.3230 1704.0400 519.8770 ;
      RECT 0.0000 518.6770 1704.3000 519.3230 ;
      RECT 0.2600 518.1230 1704.0400 518.6770 ;
      RECT 0.0000 517.4770 1704.3000 518.1230 ;
      RECT 0.2600 516.9230 1704.0400 517.4770 ;
      RECT 0.0000 516.2770 1704.3000 516.9230 ;
      RECT 0.2600 515.7230 1704.0400 516.2770 ;
      RECT 0.0000 515.0770 1704.3000 515.7230 ;
      RECT 0.2600 514.5230 1704.0400 515.0770 ;
      RECT 0.0000 513.8770 1704.3000 514.5230 ;
      RECT 0.2600 513.3230 1704.0400 513.8770 ;
      RECT 0.0000 512.6770 1704.3000 513.3230 ;
      RECT 0.2600 512.1230 1704.0400 512.6770 ;
      RECT 0.0000 511.4770 1704.3000 512.1230 ;
      RECT 0.2600 510.9230 1704.0400 511.4770 ;
      RECT 0.0000 510.2770 1704.3000 510.9230 ;
      RECT 0.2600 509.7230 1704.0400 510.2770 ;
      RECT 0.0000 509.0770 1704.3000 509.7230 ;
      RECT 0.2600 508.5230 1704.0400 509.0770 ;
      RECT 0.0000 507.8770 1704.3000 508.5230 ;
      RECT 0.2600 507.3230 1704.0400 507.8770 ;
      RECT 0.0000 506.6770 1704.3000 507.3230 ;
      RECT 0.2600 506.1230 1704.0400 506.6770 ;
      RECT 0.0000 505.4770 1704.3000 506.1230 ;
      RECT 0.2600 504.9230 1704.0400 505.4770 ;
      RECT 0.0000 504.2770 1704.3000 504.9230 ;
      RECT 0.2600 503.7230 1704.0400 504.2770 ;
      RECT 0.0000 503.0770 1704.3000 503.7230 ;
      RECT 0.2600 502.5230 1704.0400 503.0770 ;
      RECT 0.0000 501.8770 1704.3000 502.5230 ;
      RECT 0.2600 501.3230 1704.0400 501.8770 ;
      RECT 0.0000 500.6770 1704.3000 501.3230 ;
      RECT 0.2600 500.1230 1704.0400 500.6770 ;
      RECT 0.0000 499.4770 1704.3000 500.1230 ;
      RECT 0.2600 498.9230 1704.0400 499.4770 ;
      RECT 0.0000 498.2770 1704.3000 498.9230 ;
      RECT 0.2600 497.7230 1704.0400 498.2770 ;
      RECT 0.0000 497.0770 1704.3000 497.7230 ;
      RECT 0.2600 496.5230 1704.0400 497.0770 ;
      RECT 0.0000 495.8770 1704.3000 496.5230 ;
      RECT 0.2600 495.3230 1704.0400 495.8770 ;
      RECT 0.0000 494.6770 1704.3000 495.3230 ;
      RECT 0.2600 494.1230 1704.0400 494.6770 ;
      RECT 0.0000 493.4770 1704.3000 494.1230 ;
      RECT 0.2600 492.9230 1704.0400 493.4770 ;
      RECT 0.0000 492.2770 1704.3000 492.9230 ;
      RECT 0.2600 491.7230 1704.0400 492.2770 ;
      RECT 0.0000 491.0770 1704.3000 491.7230 ;
      RECT 0.2600 490.5230 1704.0400 491.0770 ;
      RECT 0.0000 489.8770 1704.3000 490.5230 ;
      RECT 0.2600 489.3230 1704.0400 489.8770 ;
      RECT 0.0000 488.6770 1704.3000 489.3230 ;
      RECT 0.2600 488.1230 1704.0400 488.6770 ;
      RECT 0.0000 487.4770 1704.3000 488.1230 ;
      RECT 0.2600 486.9230 1704.0400 487.4770 ;
      RECT 0.0000 486.2770 1704.3000 486.9230 ;
      RECT 0.2600 485.7230 1704.0400 486.2770 ;
      RECT 0.0000 485.0770 1704.3000 485.7230 ;
      RECT 0.2600 484.5230 1704.0400 485.0770 ;
      RECT 0.0000 483.8770 1704.3000 484.5230 ;
      RECT 0.2600 483.3230 1704.0400 483.8770 ;
      RECT 0.0000 482.6770 1704.3000 483.3230 ;
      RECT 0.2600 482.1230 1704.0400 482.6770 ;
      RECT 0.0000 481.4770 1704.3000 482.1230 ;
      RECT 0.2600 480.9230 1704.0400 481.4770 ;
      RECT 0.0000 480.2770 1704.3000 480.9230 ;
      RECT 0.2600 479.7230 1704.0400 480.2770 ;
      RECT 0.0000 479.0770 1704.3000 479.7230 ;
      RECT 0.2600 478.5230 1704.0400 479.0770 ;
      RECT 0.0000 477.8770 1704.3000 478.5230 ;
      RECT 0.2600 477.3230 1704.0400 477.8770 ;
      RECT 0.0000 476.6770 1704.3000 477.3230 ;
      RECT 0.2600 476.1230 1704.0400 476.6770 ;
      RECT 0.0000 475.4770 1704.3000 476.1230 ;
      RECT 0.2600 474.9230 1704.0400 475.4770 ;
      RECT 0.0000 474.2770 1704.3000 474.9230 ;
      RECT 0.2600 473.7230 1704.0400 474.2770 ;
      RECT 0.0000 473.0770 1704.3000 473.7230 ;
      RECT 0.2600 472.5230 1704.0400 473.0770 ;
      RECT 0.0000 471.8770 1704.3000 472.5230 ;
      RECT 0.2600 471.3230 1704.0400 471.8770 ;
      RECT 0.0000 470.6770 1704.3000 471.3230 ;
      RECT 0.2600 470.1230 1704.0400 470.6770 ;
      RECT 0.0000 469.4770 1704.3000 470.1230 ;
      RECT 0.2600 468.9230 1704.0400 469.4770 ;
      RECT 0.0000 468.2770 1704.3000 468.9230 ;
      RECT 0.2600 467.7230 1704.0400 468.2770 ;
      RECT 0.0000 467.0770 1704.3000 467.7230 ;
      RECT 0.2600 466.5230 1704.0400 467.0770 ;
      RECT 0.0000 465.8770 1704.3000 466.5230 ;
      RECT 0.2600 465.3230 1704.0400 465.8770 ;
      RECT 0.0000 464.6770 1704.3000 465.3230 ;
      RECT 0.2600 464.1230 1704.0400 464.6770 ;
      RECT 0.0000 463.4770 1704.3000 464.1230 ;
      RECT 0.2600 462.9230 1704.0400 463.4770 ;
      RECT 0.0000 462.2770 1704.3000 462.9230 ;
      RECT 0.2600 461.7230 1704.0400 462.2770 ;
      RECT 0.0000 461.0770 1704.3000 461.7230 ;
      RECT 0.2600 460.5230 1704.0400 461.0770 ;
      RECT 0.0000 459.8770 1704.3000 460.5230 ;
      RECT 0.2600 459.3230 1704.0400 459.8770 ;
      RECT 0.0000 458.6770 1704.3000 459.3230 ;
      RECT 0.2600 458.1230 1704.0400 458.6770 ;
      RECT 0.0000 457.4770 1704.3000 458.1230 ;
      RECT 0.2600 456.9230 1704.0400 457.4770 ;
      RECT 0.0000 456.2770 1704.3000 456.9230 ;
      RECT 0.2600 455.7230 1704.0400 456.2770 ;
      RECT 0.0000 455.0770 1704.3000 455.7230 ;
      RECT 0.2600 454.5230 1704.0400 455.0770 ;
      RECT 0.0000 453.8770 1704.3000 454.5230 ;
      RECT 0.2600 453.3230 1704.0400 453.8770 ;
      RECT 0.0000 452.6770 1704.3000 453.3230 ;
      RECT 0.2600 452.1230 1704.0400 452.6770 ;
      RECT 0.0000 451.4770 1704.3000 452.1230 ;
      RECT 0.2600 450.9230 1704.0400 451.4770 ;
      RECT 0.0000 450.2770 1704.3000 450.9230 ;
      RECT 0.2600 449.7230 1704.0400 450.2770 ;
      RECT 0.0000 449.0770 1704.3000 449.7230 ;
      RECT 0.2600 448.5230 1704.0400 449.0770 ;
      RECT 0.0000 447.8770 1704.3000 448.5230 ;
      RECT 0.2600 447.3230 1704.0400 447.8770 ;
      RECT 0.0000 446.6770 1704.3000 447.3230 ;
      RECT 0.2600 446.1230 1704.0400 446.6770 ;
      RECT 0.0000 445.4770 1704.3000 446.1230 ;
      RECT 0.2600 444.9230 1704.0400 445.4770 ;
      RECT 0.0000 444.2770 1704.3000 444.9230 ;
      RECT 0.2600 443.7230 1704.0400 444.2770 ;
      RECT 0.0000 443.0770 1704.3000 443.7230 ;
      RECT 0.2600 442.5230 1704.0400 443.0770 ;
      RECT 0.0000 441.8770 1704.3000 442.5230 ;
      RECT 0.2600 441.3230 1704.0400 441.8770 ;
      RECT 0.0000 440.6770 1704.3000 441.3230 ;
      RECT 0.2600 440.1230 1704.0400 440.6770 ;
      RECT 0.0000 439.4770 1704.3000 440.1230 ;
      RECT 0.2600 438.9230 1704.0400 439.4770 ;
      RECT 0.0000 438.2770 1704.3000 438.9230 ;
      RECT 0.2600 437.7230 1704.0400 438.2770 ;
      RECT 0.0000 437.0770 1704.3000 437.7230 ;
      RECT 0.2600 436.5230 1704.0400 437.0770 ;
      RECT 0.0000 435.8770 1704.3000 436.5230 ;
      RECT 0.2600 435.3230 1704.0400 435.8770 ;
      RECT 0.0000 434.6770 1704.3000 435.3230 ;
      RECT 0.2600 434.1230 1704.0400 434.6770 ;
      RECT 0.0000 433.4770 1704.3000 434.1230 ;
      RECT 0.2600 432.9230 1704.0400 433.4770 ;
      RECT 0.0000 432.2770 1704.3000 432.9230 ;
      RECT 0.2600 431.7230 1704.0400 432.2770 ;
      RECT 0.0000 431.0770 1704.3000 431.7230 ;
      RECT 0.2600 430.5230 1704.0400 431.0770 ;
      RECT 0.0000 429.8770 1704.3000 430.5230 ;
      RECT 0.2600 429.3230 1704.0400 429.8770 ;
      RECT 0.0000 428.6770 1704.3000 429.3230 ;
      RECT 0.2600 428.1230 1704.0400 428.6770 ;
      RECT 0.0000 427.4770 1704.3000 428.1230 ;
      RECT 0.2600 426.9230 1704.0400 427.4770 ;
      RECT 0.0000 426.2770 1704.3000 426.9230 ;
      RECT 0.2600 425.7230 1704.0400 426.2770 ;
      RECT 0.0000 425.0770 1704.3000 425.7230 ;
      RECT 0.2600 424.5230 1704.0400 425.0770 ;
      RECT 0.0000 423.8770 1704.3000 424.5230 ;
      RECT 0.2600 423.3230 1704.0400 423.8770 ;
      RECT 0.0000 422.6770 1704.3000 423.3230 ;
      RECT 0.2600 422.1230 1704.0400 422.6770 ;
      RECT 0.0000 421.4770 1704.3000 422.1230 ;
      RECT 0.2600 420.9230 1704.0400 421.4770 ;
      RECT 0.0000 420.2770 1704.3000 420.9230 ;
      RECT 0.2600 419.7230 1704.0400 420.2770 ;
      RECT 0.0000 419.0770 1704.3000 419.7230 ;
      RECT 0.2600 418.5230 1704.0400 419.0770 ;
      RECT 0.0000 417.8770 1704.3000 418.5230 ;
      RECT 0.2600 417.3230 1704.0400 417.8770 ;
      RECT 0.0000 416.6770 1704.3000 417.3230 ;
      RECT 0.2600 416.1230 1704.0400 416.6770 ;
      RECT 0.0000 415.4770 1704.3000 416.1230 ;
      RECT 0.2600 414.9230 1704.0400 415.4770 ;
      RECT 0.0000 414.2770 1704.3000 414.9230 ;
      RECT 0.2600 413.7230 1704.0400 414.2770 ;
      RECT 0.0000 413.0770 1704.3000 413.7230 ;
      RECT 0.2600 412.5230 1704.0400 413.0770 ;
      RECT 0.0000 411.8770 1704.3000 412.5230 ;
      RECT 0.2600 411.3230 1704.0400 411.8770 ;
      RECT 0.0000 410.6770 1704.3000 411.3230 ;
      RECT 0.2600 410.1230 1704.0400 410.6770 ;
      RECT 0.0000 409.4770 1704.3000 410.1230 ;
      RECT 0.2600 408.9230 1704.0400 409.4770 ;
      RECT 0.0000 408.2770 1704.3000 408.9230 ;
      RECT 0.2600 407.7230 1704.0400 408.2770 ;
      RECT 0.0000 407.0770 1704.3000 407.7230 ;
      RECT 0.2600 406.5230 1704.0400 407.0770 ;
      RECT 0.0000 405.8770 1704.3000 406.5230 ;
      RECT 0.2600 405.3230 1704.0400 405.8770 ;
      RECT 0.0000 404.6770 1704.3000 405.3230 ;
      RECT 0.2600 404.1230 1704.0400 404.6770 ;
      RECT 0.0000 403.4770 1704.3000 404.1230 ;
      RECT 0.2600 402.9230 1704.0400 403.4770 ;
      RECT 0.0000 402.2770 1704.3000 402.9230 ;
      RECT 0.2600 401.7230 1704.0400 402.2770 ;
      RECT 0.0000 401.0770 1704.3000 401.7230 ;
      RECT 0.2600 400.5230 1704.0400 401.0770 ;
      RECT 0.0000 399.8770 1704.3000 400.5230 ;
      RECT 0.2600 399.3230 1704.0400 399.8770 ;
      RECT 0.0000 398.6770 1704.3000 399.3230 ;
      RECT 0.2600 398.1230 1704.0400 398.6770 ;
      RECT 0.0000 397.4770 1704.3000 398.1230 ;
      RECT 0.2600 396.9230 1704.0400 397.4770 ;
      RECT 0.0000 396.2770 1704.3000 396.9230 ;
      RECT 0.2600 395.7230 1704.0400 396.2770 ;
      RECT 0.0000 395.0770 1704.3000 395.7230 ;
      RECT 0.2600 394.5230 1704.0400 395.0770 ;
      RECT 0.0000 393.8770 1704.3000 394.5230 ;
      RECT 0.2600 393.3230 1704.0400 393.8770 ;
      RECT 0.0000 392.6770 1704.3000 393.3230 ;
      RECT 0.2600 392.1230 1704.0400 392.6770 ;
      RECT 0.0000 391.4770 1704.3000 392.1230 ;
      RECT 0.2600 390.9230 1704.0400 391.4770 ;
      RECT 0.0000 390.2770 1704.3000 390.9230 ;
      RECT 0.2600 389.7230 1704.0400 390.2770 ;
      RECT 0.0000 389.0770 1704.3000 389.7230 ;
      RECT 0.2600 388.5230 1704.0400 389.0770 ;
      RECT 0.0000 387.8770 1704.3000 388.5230 ;
      RECT 0.2600 387.3230 1704.0400 387.8770 ;
      RECT 0.0000 386.6770 1704.3000 387.3230 ;
      RECT 0.2600 386.1230 1704.0400 386.6770 ;
      RECT 0.0000 385.4770 1704.3000 386.1230 ;
      RECT 0.2600 384.9230 1704.0400 385.4770 ;
      RECT 0.0000 384.2770 1704.3000 384.9230 ;
      RECT 0.2600 383.7230 1704.0400 384.2770 ;
      RECT 0.0000 383.0770 1704.3000 383.7230 ;
      RECT 0.2600 382.5230 1704.0400 383.0770 ;
      RECT 0.0000 381.8770 1704.3000 382.5230 ;
      RECT 0.2600 381.3230 1704.0400 381.8770 ;
      RECT 0.0000 380.6770 1704.3000 381.3230 ;
      RECT 0.2600 380.1230 1704.0400 380.6770 ;
      RECT 0.0000 379.4770 1704.3000 380.1230 ;
      RECT 0.2600 378.9230 1704.0400 379.4770 ;
      RECT 0.0000 378.2770 1704.3000 378.9230 ;
      RECT 0.2600 377.7230 1704.0400 378.2770 ;
      RECT 0.0000 377.0770 1704.3000 377.7230 ;
      RECT 0.2600 376.5230 1704.0400 377.0770 ;
      RECT 0.0000 375.8770 1704.3000 376.5230 ;
      RECT 0.2600 375.3230 1704.0400 375.8770 ;
      RECT 0.0000 374.6770 1704.3000 375.3230 ;
      RECT 0.2600 374.1230 1704.0400 374.6770 ;
      RECT 0.0000 373.4770 1704.3000 374.1230 ;
      RECT 0.2600 372.9230 1704.0400 373.4770 ;
      RECT 0.0000 372.2770 1704.3000 372.9230 ;
      RECT 0.2600 371.7230 1704.0400 372.2770 ;
      RECT 0.0000 371.0770 1704.3000 371.7230 ;
      RECT 0.2600 370.5230 1704.0400 371.0770 ;
      RECT 0.0000 369.8770 1704.3000 370.5230 ;
      RECT 0.2600 369.3230 1704.0400 369.8770 ;
      RECT 0.0000 368.6770 1704.3000 369.3230 ;
      RECT 0.2600 368.1230 1704.0400 368.6770 ;
      RECT 0.0000 367.4770 1704.3000 368.1230 ;
      RECT 0.2600 366.9230 1704.0400 367.4770 ;
      RECT 0.0000 366.2770 1704.3000 366.9230 ;
      RECT 0.2600 365.7230 1704.0400 366.2770 ;
      RECT 0.0000 365.0770 1704.3000 365.7230 ;
      RECT 0.2600 364.5230 1704.0400 365.0770 ;
      RECT 0.0000 363.8770 1704.3000 364.5230 ;
      RECT 0.2600 363.3230 1704.0400 363.8770 ;
      RECT 0.0000 362.6770 1704.3000 363.3230 ;
      RECT 0.2600 362.1230 1704.0400 362.6770 ;
      RECT 0.0000 361.4770 1704.3000 362.1230 ;
      RECT 0.2600 360.9230 1704.0400 361.4770 ;
      RECT 0.0000 360.2770 1704.3000 360.9230 ;
      RECT 0.2600 359.7230 1704.0400 360.2770 ;
      RECT 0.0000 359.0770 1704.3000 359.7230 ;
      RECT 0.2600 358.5230 1704.0400 359.0770 ;
      RECT 0.0000 357.8770 1704.3000 358.5230 ;
      RECT 0.2600 357.3230 1704.0400 357.8770 ;
      RECT 0.0000 356.6770 1704.3000 357.3230 ;
      RECT 0.2600 356.1230 1704.0400 356.6770 ;
      RECT 0.0000 355.4770 1704.3000 356.1230 ;
      RECT 0.2600 354.9230 1704.0400 355.4770 ;
      RECT 0.0000 354.2770 1704.3000 354.9230 ;
      RECT 0.2600 353.7230 1704.0400 354.2770 ;
      RECT 0.0000 353.0770 1704.3000 353.7230 ;
      RECT 0.2600 352.5230 1704.0400 353.0770 ;
      RECT 0.0000 351.8770 1704.3000 352.5230 ;
      RECT 0.2600 351.3230 1704.0400 351.8770 ;
      RECT 0.0000 350.6770 1704.3000 351.3230 ;
      RECT 0.2600 350.1230 1704.0400 350.6770 ;
      RECT 0.0000 349.4770 1704.3000 350.1230 ;
      RECT 0.2600 348.9230 1704.0400 349.4770 ;
      RECT 0.0000 348.2770 1704.3000 348.9230 ;
      RECT 0.2600 347.7230 1704.0400 348.2770 ;
      RECT 0.0000 347.0770 1704.3000 347.7230 ;
      RECT 0.2600 346.5230 1704.0400 347.0770 ;
      RECT 0.0000 345.8770 1704.3000 346.5230 ;
      RECT 0.2600 345.3230 1704.0400 345.8770 ;
      RECT 0.0000 344.6770 1704.3000 345.3230 ;
      RECT 0.2600 344.1230 1704.0400 344.6770 ;
      RECT 0.0000 343.4770 1704.3000 344.1230 ;
      RECT 0.2600 342.9230 1704.0400 343.4770 ;
      RECT 0.0000 342.2770 1704.3000 342.9230 ;
      RECT 0.2600 341.7230 1704.0400 342.2770 ;
      RECT 0.0000 341.0770 1704.3000 341.7230 ;
      RECT 0.2600 340.5230 1704.0400 341.0770 ;
      RECT 0.0000 339.8770 1704.3000 340.5230 ;
      RECT 0.2600 339.3230 1704.0400 339.8770 ;
      RECT 0.0000 338.6770 1704.3000 339.3230 ;
      RECT 0.2600 338.1230 1704.0400 338.6770 ;
      RECT 0.0000 337.4770 1704.3000 338.1230 ;
      RECT 0.2600 336.9230 1704.0400 337.4770 ;
      RECT 0.0000 336.2770 1704.3000 336.9230 ;
      RECT 0.2600 335.7230 1704.0400 336.2770 ;
      RECT 0.0000 335.0770 1704.3000 335.7230 ;
      RECT 0.2600 334.5230 1704.0400 335.0770 ;
      RECT 0.0000 333.8770 1704.3000 334.5230 ;
      RECT 0.2600 333.3230 1704.0400 333.8770 ;
      RECT 0.0000 332.6770 1704.3000 333.3230 ;
      RECT 0.2600 332.1230 1704.0400 332.6770 ;
      RECT 0.0000 331.4770 1704.3000 332.1230 ;
      RECT 0.2600 330.9230 1704.0400 331.4770 ;
      RECT 0.0000 330.2770 1704.3000 330.9230 ;
      RECT 0.2600 329.7230 1704.0400 330.2770 ;
      RECT 0.0000 329.0770 1704.3000 329.7230 ;
      RECT 0.2600 328.5230 1704.0400 329.0770 ;
      RECT 0.0000 327.8770 1704.3000 328.5230 ;
      RECT 0.2600 327.3230 1704.0400 327.8770 ;
      RECT 0.0000 326.6770 1704.3000 327.3230 ;
      RECT 0.2600 326.1230 1704.0400 326.6770 ;
      RECT 0.0000 325.4770 1704.3000 326.1230 ;
      RECT 0.2600 324.9230 1704.0400 325.4770 ;
      RECT 0.0000 324.2770 1704.3000 324.9230 ;
      RECT 0.2600 323.7230 1704.0400 324.2770 ;
      RECT 0.0000 323.0770 1704.3000 323.7230 ;
      RECT 0.2600 322.5230 1704.0400 323.0770 ;
      RECT 0.0000 321.8770 1704.3000 322.5230 ;
      RECT 0.2600 321.3230 1704.0400 321.8770 ;
      RECT 0.0000 320.6770 1704.3000 321.3230 ;
      RECT 0.2600 320.1230 1704.0400 320.6770 ;
      RECT 0.0000 319.4770 1704.3000 320.1230 ;
      RECT 0.2600 318.9230 1704.0400 319.4770 ;
      RECT 0.0000 318.2770 1704.3000 318.9230 ;
      RECT 0.2600 317.7230 1704.0400 318.2770 ;
      RECT 0.0000 317.0770 1704.3000 317.7230 ;
      RECT 0.2600 316.5230 1704.0400 317.0770 ;
      RECT 0.0000 315.8770 1704.3000 316.5230 ;
      RECT 0.2600 315.3230 1704.0400 315.8770 ;
      RECT 0.0000 314.6770 1704.3000 315.3230 ;
      RECT 0.2600 314.1230 1704.0400 314.6770 ;
      RECT 0.0000 313.4770 1704.3000 314.1230 ;
      RECT 0.2600 312.9230 1704.0400 313.4770 ;
      RECT 0.0000 312.2770 1704.3000 312.9230 ;
      RECT 0.2600 311.7230 1704.0400 312.2770 ;
      RECT 0.0000 311.0770 1704.3000 311.7230 ;
      RECT 0.2600 310.5230 1704.0400 311.0770 ;
      RECT 0.0000 309.8770 1704.3000 310.5230 ;
      RECT 0.2600 309.3230 1704.0400 309.8770 ;
      RECT 0.0000 308.6770 1704.3000 309.3230 ;
      RECT 0.2600 308.1230 1704.0400 308.6770 ;
      RECT 0.0000 307.4770 1704.3000 308.1230 ;
      RECT 0.2600 306.9230 1704.0400 307.4770 ;
      RECT 0.0000 306.2770 1704.3000 306.9230 ;
      RECT 0.2600 305.7230 1704.0400 306.2770 ;
      RECT 0.0000 305.0770 1704.3000 305.7230 ;
      RECT 0.2600 304.5230 1704.0400 305.0770 ;
      RECT 0.0000 303.8770 1704.3000 304.5230 ;
      RECT 0.2600 303.3230 1704.0400 303.8770 ;
      RECT 0.0000 302.6770 1704.3000 303.3230 ;
      RECT 0.2600 302.1230 1704.0400 302.6770 ;
      RECT 0.0000 301.4770 1704.3000 302.1230 ;
      RECT 0.2600 300.9230 1704.0400 301.4770 ;
      RECT 0.0000 300.2770 1704.3000 300.9230 ;
      RECT 0.2600 299.7230 1704.0400 300.2770 ;
      RECT 0.0000 299.0770 1704.3000 299.7230 ;
      RECT 0.2600 298.5230 1704.0400 299.0770 ;
      RECT 0.0000 297.8770 1704.3000 298.5230 ;
      RECT 0.2600 297.3230 1704.0400 297.8770 ;
      RECT 0.0000 296.6770 1704.3000 297.3230 ;
      RECT 0.2600 296.1230 1704.0400 296.6770 ;
      RECT 0.0000 295.4770 1704.3000 296.1230 ;
      RECT 0.2600 294.9230 1704.0400 295.4770 ;
      RECT 0.0000 294.2770 1704.3000 294.9230 ;
      RECT 0.2600 293.7230 1704.0400 294.2770 ;
      RECT 0.0000 293.0770 1704.3000 293.7230 ;
      RECT 0.2600 292.5230 1704.0400 293.0770 ;
      RECT 0.0000 291.8770 1704.3000 292.5230 ;
      RECT 0.2600 291.3230 1704.0400 291.8770 ;
      RECT 0.0000 290.6770 1704.3000 291.3230 ;
      RECT 0.2600 290.1230 1704.0400 290.6770 ;
      RECT 0.0000 289.4770 1704.3000 290.1230 ;
      RECT 0.2600 288.9230 1704.0400 289.4770 ;
      RECT 0.0000 288.2770 1704.3000 288.9230 ;
      RECT 0.2600 287.7230 1704.0400 288.2770 ;
      RECT 0.0000 287.0770 1704.3000 287.7230 ;
      RECT 0.2600 286.5230 1704.0400 287.0770 ;
      RECT 0.0000 285.8770 1704.3000 286.5230 ;
      RECT 0.2600 285.3230 1704.0400 285.8770 ;
      RECT 0.0000 284.6770 1704.3000 285.3230 ;
      RECT 0.2600 284.1230 1704.0400 284.6770 ;
      RECT 0.0000 283.4770 1704.3000 284.1230 ;
      RECT 0.2600 282.9230 1704.0400 283.4770 ;
      RECT 0.0000 282.2770 1704.3000 282.9230 ;
      RECT 0.2600 281.7230 1704.0400 282.2770 ;
      RECT 0.0000 281.0770 1704.3000 281.7230 ;
      RECT 0.2600 280.5230 1704.0400 281.0770 ;
      RECT 0.0000 279.8770 1704.3000 280.5230 ;
      RECT 0.2600 279.3230 1704.0400 279.8770 ;
      RECT 0.0000 278.6770 1704.3000 279.3230 ;
      RECT 0.2600 278.1230 1704.0400 278.6770 ;
      RECT 0.0000 277.4770 1704.3000 278.1230 ;
      RECT 0.2600 276.9230 1704.0400 277.4770 ;
      RECT 0.0000 276.2770 1704.3000 276.9230 ;
      RECT 0.2600 275.7230 1704.0400 276.2770 ;
      RECT 0.0000 275.0770 1704.3000 275.7230 ;
      RECT 0.2600 274.5230 1704.0400 275.0770 ;
      RECT 0.0000 273.8770 1704.3000 274.5230 ;
      RECT 0.2600 273.3230 1704.0400 273.8770 ;
      RECT 0.0000 272.6770 1704.3000 273.3230 ;
      RECT 0.2600 272.1230 1704.0400 272.6770 ;
      RECT 0.0000 271.4770 1704.3000 272.1230 ;
      RECT 0.2600 270.9230 1704.0400 271.4770 ;
      RECT 0.0000 270.2770 1704.3000 270.9230 ;
      RECT 0.2600 269.7230 1704.0400 270.2770 ;
      RECT 0.0000 269.0770 1704.3000 269.7230 ;
      RECT 0.2600 268.5230 1704.0400 269.0770 ;
      RECT 0.0000 267.8770 1704.3000 268.5230 ;
      RECT 0.2600 267.3230 1704.0400 267.8770 ;
      RECT 0.0000 266.6770 1704.3000 267.3230 ;
      RECT 0.2600 266.1230 1704.0400 266.6770 ;
      RECT 0.0000 265.4770 1704.3000 266.1230 ;
      RECT 0.2600 264.9230 1704.0400 265.4770 ;
      RECT 0.0000 264.2770 1704.3000 264.9230 ;
      RECT 0.2600 263.7230 1704.0400 264.2770 ;
      RECT 0.0000 263.0770 1704.3000 263.7230 ;
      RECT 0.2600 262.5230 1704.0400 263.0770 ;
      RECT 0.0000 261.8770 1704.3000 262.5230 ;
      RECT 0.2600 261.3230 1704.0400 261.8770 ;
      RECT 0.0000 260.6770 1704.3000 261.3230 ;
      RECT 0.2600 260.1230 1704.0400 260.6770 ;
      RECT 0.0000 259.4770 1704.3000 260.1230 ;
      RECT 0.2600 258.9230 1704.0400 259.4770 ;
      RECT 0.0000 258.2770 1704.3000 258.9230 ;
      RECT 0.2600 257.7230 1704.0400 258.2770 ;
      RECT 0.0000 257.0770 1704.3000 257.7230 ;
      RECT 0.2600 256.5230 1704.0400 257.0770 ;
      RECT 0.0000 255.8770 1704.3000 256.5230 ;
      RECT 0.2600 255.3230 1704.0400 255.8770 ;
      RECT 0.0000 254.6770 1704.3000 255.3230 ;
      RECT 0.2600 254.1230 1704.0400 254.6770 ;
      RECT 0.0000 253.4770 1704.3000 254.1230 ;
      RECT 0.2600 252.9230 1704.0400 253.4770 ;
      RECT 0.0000 252.2770 1704.3000 252.9230 ;
      RECT 0.2600 251.7230 1704.0400 252.2770 ;
      RECT 0.0000 251.0770 1704.3000 251.7230 ;
      RECT 0.2600 250.5230 1704.0400 251.0770 ;
      RECT 0.0000 249.8770 1704.3000 250.5230 ;
      RECT 0.2600 249.3230 1704.0400 249.8770 ;
      RECT 0.0000 248.6770 1704.3000 249.3230 ;
      RECT 0.2600 248.1230 1704.0400 248.6770 ;
      RECT 0.0000 247.4770 1704.3000 248.1230 ;
      RECT 0.2600 246.9230 1704.0400 247.4770 ;
      RECT 0.0000 246.2770 1704.3000 246.9230 ;
      RECT 0.2600 245.7230 1704.0400 246.2770 ;
      RECT 0.0000 245.0770 1704.3000 245.7230 ;
      RECT 0.2600 244.5230 1704.0400 245.0770 ;
      RECT 0.0000 243.8770 1704.3000 244.5230 ;
      RECT 0.2600 243.3230 1704.0400 243.8770 ;
      RECT 0.0000 242.6770 1704.3000 243.3230 ;
      RECT 0.2600 242.1230 1704.0400 242.6770 ;
      RECT 0.0000 241.4770 1704.3000 242.1230 ;
      RECT 0.2600 240.9230 1704.0400 241.4770 ;
      RECT 0.0000 240.2770 1704.3000 240.9230 ;
      RECT 0.2600 239.7230 1704.0400 240.2770 ;
      RECT 0.0000 239.0770 1704.3000 239.7230 ;
      RECT 0.2600 238.5230 1704.0400 239.0770 ;
      RECT 0.0000 237.8770 1704.3000 238.5230 ;
      RECT 0.2600 237.3230 1704.0400 237.8770 ;
      RECT 0.0000 236.6770 1704.3000 237.3230 ;
      RECT 0.2600 236.1230 1704.0400 236.6770 ;
      RECT 0.0000 235.4770 1704.3000 236.1230 ;
      RECT 0.2600 234.9230 1704.0400 235.4770 ;
      RECT 0.0000 234.2770 1704.3000 234.9230 ;
      RECT 0.2600 233.7230 1704.0400 234.2770 ;
      RECT 0.0000 233.0770 1704.3000 233.7230 ;
      RECT 0.2600 232.5230 1704.0400 233.0770 ;
      RECT 0.0000 231.8770 1704.3000 232.5230 ;
      RECT 0.2600 231.3230 1704.0400 231.8770 ;
      RECT 0.0000 230.6770 1704.3000 231.3230 ;
      RECT 0.2600 230.1230 1704.0400 230.6770 ;
      RECT 0.0000 229.4770 1704.3000 230.1230 ;
      RECT 0.2600 228.9230 1704.0400 229.4770 ;
      RECT 0.0000 228.2770 1704.3000 228.9230 ;
      RECT 0.2600 227.7230 1704.0400 228.2770 ;
      RECT 0.0000 227.0770 1704.3000 227.7230 ;
      RECT 0.2600 226.5230 1704.0400 227.0770 ;
      RECT 0.0000 225.8770 1704.3000 226.5230 ;
      RECT 0.2600 225.3230 1704.0400 225.8770 ;
      RECT 0.0000 224.6770 1704.3000 225.3230 ;
      RECT 0.2600 224.1230 1704.0400 224.6770 ;
      RECT 0.0000 223.4770 1704.3000 224.1230 ;
      RECT 0.2600 222.9230 1704.0400 223.4770 ;
      RECT 0.0000 222.2770 1704.3000 222.9230 ;
      RECT 0.2600 221.7230 1704.0400 222.2770 ;
      RECT 0.0000 221.0770 1704.3000 221.7230 ;
      RECT 0.2600 220.5230 1704.0400 221.0770 ;
      RECT 0.0000 219.8770 1704.3000 220.5230 ;
      RECT 0.2600 219.3230 1704.0400 219.8770 ;
      RECT 0.0000 218.6770 1704.3000 219.3230 ;
      RECT 0.2600 218.1230 1704.0400 218.6770 ;
      RECT 0.0000 217.4770 1704.3000 218.1230 ;
      RECT 0.2600 216.9230 1704.0400 217.4770 ;
      RECT 0.0000 216.2770 1704.3000 216.9230 ;
      RECT 0.2600 215.7230 1704.0400 216.2770 ;
      RECT 0.0000 215.0770 1704.3000 215.7230 ;
      RECT 0.2600 214.5230 1704.0400 215.0770 ;
      RECT 0.0000 213.8770 1704.3000 214.5230 ;
      RECT 0.2600 213.3230 1704.0400 213.8770 ;
      RECT 0.0000 212.6770 1704.3000 213.3230 ;
      RECT 0.2600 212.1230 1704.0400 212.6770 ;
      RECT 0.0000 211.4770 1704.3000 212.1230 ;
      RECT 0.2600 210.9230 1704.0400 211.4770 ;
      RECT 0.0000 210.2770 1704.3000 210.9230 ;
      RECT 0.2600 209.7230 1704.0400 210.2770 ;
      RECT 0.0000 209.0770 1704.3000 209.7230 ;
      RECT 0.2600 208.5230 1704.0400 209.0770 ;
      RECT 0.0000 207.8770 1704.3000 208.5230 ;
      RECT 0.2600 207.3230 1704.0400 207.8770 ;
      RECT 0.0000 206.6770 1704.3000 207.3230 ;
      RECT 0.2600 206.1230 1704.0400 206.6770 ;
      RECT 0.0000 205.4770 1704.3000 206.1230 ;
      RECT 0.2600 204.9230 1704.0400 205.4770 ;
      RECT 0.0000 204.2770 1704.3000 204.9230 ;
      RECT 0.2600 203.7230 1704.0400 204.2770 ;
      RECT 0.0000 203.0770 1704.3000 203.7230 ;
      RECT 0.2600 202.5230 1704.0400 203.0770 ;
      RECT 0.0000 201.8770 1704.3000 202.5230 ;
      RECT 0.2600 201.3230 1704.0400 201.8770 ;
      RECT 0.0000 200.6770 1704.3000 201.3230 ;
      RECT 0.2600 200.1230 1704.0400 200.6770 ;
      RECT 0.0000 199.4770 1704.3000 200.1230 ;
      RECT 0.2600 198.9230 1704.0400 199.4770 ;
      RECT 0.0000 198.2770 1704.3000 198.9230 ;
      RECT 0.2600 197.7230 1704.0400 198.2770 ;
      RECT 0.0000 197.0770 1704.3000 197.7230 ;
      RECT 0.2600 196.5230 1704.0400 197.0770 ;
      RECT 0.0000 195.8770 1704.3000 196.5230 ;
      RECT 0.2600 195.3230 1704.0400 195.8770 ;
      RECT 0.0000 194.6770 1704.3000 195.3230 ;
      RECT 0.2600 194.1230 1704.0400 194.6770 ;
      RECT 0.0000 193.4770 1704.3000 194.1230 ;
      RECT 0.2600 192.9230 1704.0400 193.4770 ;
      RECT 0.0000 192.2770 1704.3000 192.9230 ;
      RECT 0.2600 191.7230 1704.0400 192.2770 ;
      RECT 0.0000 191.0770 1704.3000 191.7230 ;
      RECT 0.2600 190.5230 1704.0400 191.0770 ;
      RECT 0.0000 189.8770 1704.3000 190.5230 ;
      RECT 0.2600 189.3230 1704.0400 189.8770 ;
      RECT 0.0000 188.6770 1704.3000 189.3230 ;
      RECT 0.2600 188.1230 1704.0400 188.6770 ;
      RECT 0.0000 187.4770 1704.3000 188.1230 ;
      RECT 0.2600 186.9230 1704.0400 187.4770 ;
      RECT 0.0000 186.2770 1704.3000 186.9230 ;
      RECT 0.2600 185.7230 1704.0400 186.2770 ;
      RECT 0.0000 185.0770 1704.3000 185.7230 ;
      RECT 0.2600 184.5230 1704.0400 185.0770 ;
      RECT 0.0000 183.8770 1704.3000 184.5230 ;
      RECT 0.2600 183.3230 1704.0400 183.8770 ;
      RECT 0.0000 182.6770 1704.3000 183.3230 ;
      RECT 0.2600 182.1230 1704.0400 182.6770 ;
      RECT 0.0000 181.4770 1704.3000 182.1230 ;
      RECT 0.2600 180.9230 1704.0400 181.4770 ;
      RECT 0.0000 180.2770 1704.3000 180.9230 ;
      RECT 0.2600 179.7230 1704.0400 180.2770 ;
      RECT 0.0000 179.0770 1704.3000 179.7230 ;
      RECT 0.2600 178.5230 1704.0400 179.0770 ;
      RECT 0.0000 177.8770 1704.3000 178.5230 ;
      RECT 0.2600 177.3230 1704.0400 177.8770 ;
      RECT 0.0000 176.6770 1704.3000 177.3230 ;
      RECT 0.2600 176.1230 1704.0400 176.6770 ;
      RECT 0.0000 175.4770 1704.3000 176.1230 ;
      RECT 0.2600 174.9230 1704.0400 175.4770 ;
      RECT 0.0000 174.2770 1704.3000 174.9230 ;
      RECT 0.2600 173.7230 1704.0400 174.2770 ;
      RECT 0.0000 173.0770 1704.3000 173.7230 ;
      RECT 0.2600 172.5230 1704.0400 173.0770 ;
      RECT 0.0000 171.8770 1704.3000 172.5230 ;
      RECT 0.2600 171.3230 1704.0400 171.8770 ;
      RECT 0.0000 170.6770 1704.3000 171.3230 ;
      RECT 0.2600 170.1230 1704.0400 170.6770 ;
      RECT 0.0000 169.4770 1704.3000 170.1230 ;
      RECT 0.2600 168.9230 1704.0400 169.4770 ;
      RECT 0.0000 168.2770 1704.3000 168.9230 ;
      RECT 0.2600 167.7230 1704.0400 168.2770 ;
      RECT 0.0000 167.0770 1704.3000 167.7230 ;
      RECT 0.2600 166.5230 1704.0400 167.0770 ;
      RECT 0.0000 165.8770 1704.3000 166.5230 ;
      RECT 0.2600 165.3230 1704.0400 165.8770 ;
      RECT 0.0000 164.6770 1704.3000 165.3230 ;
      RECT 0.2600 164.1230 1704.0400 164.6770 ;
      RECT 0.0000 163.4770 1704.3000 164.1230 ;
      RECT 0.2600 162.9230 1704.0400 163.4770 ;
      RECT 0.0000 162.2770 1704.3000 162.9230 ;
      RECT 0.2600 161.7230 1704.0400 162.2770 ;
      RECT 0.0000 161.0770 1704.3000 161.7230 ;
      RECT 0.2600 160.5230 1704.0400 161.0770 ;
      RECT 0.0000 159.8770 1704.3000 160.5230 ;
      RECT 0.2600 159.3230 1704.0400 159.8770 ;
      RECT 0.0000 158.6770 1704.3000 159.3230 ;
      RECT 0.2600 158.1230 1704.0400 158.6770 ;
      RECT 0.0000 157.4770 1704.3000 158.1230 ;
      RECT 0.2600 156.9230 1704.0400 157.4770 ;
      RECT 0.0000 156.2770 1704.3000 156.9230 ;
      RECT 0.2600 155.7230 1704.0400 156.2770 ;
      RECT 0.0000 155.0770 1704.3000 155.7230 ;
      RECT 0.2600 154.5230 1704.0400 155.0770 ;
      RECT 0.0000 153.8770 1704.3000 154.5230 ;
      RECT 0.2600 153.3230 1704.0400 153.8770 ;
      RECT 0.0000 152.6770 1704.3000 153.3230 ;
      RECT 0.2600 152.1230 1704.0400 152.6770 ;
      RECT 0.0000 151.4770 1704.3000 152.1230 ;
      RECT 0.2600 150.9230 1704.0400 151.4770 ;
      RECT 0.0000 150.2770 1704.3000 150.9230 ;
      RECT 0.2600 149.7230 1704.0400 150.2770 ;
      RECT 0.0000 149.0770 1704.3000 149.7230 ;
      RECT 0.2600 148.5230 1704.0400 149.0770 ;
      RECT 0.0000 147.8770 1704.3000 148.5230 ;
      RECT 0.2600 147.3230 1704.0400 147.8770 ;
      RECT 0.0000 146.6770 1704.3000 147.3230 ;
      RECT 0.2600 146.1230 1704.0400 146.6770 ;
      RECT 0.0000 145.4770 1704.3000 146.1230 ;
      RECT 0.2600 144.9230 1704.0400 145.4770 ;
      RECT 0.0000 144.2770 1704.3000 144.9230 ;
      RECT 0.2600 143.7230 1704.0400 144.2770 ;
      RECT 0.0000 143.0770 1704.3000 143.7230 ;
      RECT 0.2600 142.5230 1704.0400 143.0770 ;
      RECT 0.0000 141.8770 1704.3000 142.5230 ;
      RECT 0.2600 141.3230 1704.0400 141.8770 ;
      RECT 0.0000 140.6770 1704.3000 141.3230 ;
      RECT 0.2600 140.1230 1704.0400 140.6770 ;
      RECT 0.0000 139.4770 1704.3000 140.1230 ;
      RECT 0.2600 138.9230 1704.0400 139.4770 ;
      RECT 0.0000 138.2770 1704.3000 138.9230 ;
      RECT 0.2600 137.7230 1704.0400 138.2770 ;
      RECT 0.0000 137.0770 1704.3000 137.7230 ;
      RECT 0.2600 136.5230 1704.0400 137.0770 ;
      RECT 0.0000 135.8770 1704.3000 136.5230 ;
      RECT 0.2600 135.3230 1704.0400 135.8770 ;
      RECT 0.0000 134.6770 1704.3000 135.3230 ;
      RECT 0.2600 134.1230 1704.0400 134.6770 ;
      RECT 0.0000 133.4770 1704.3000 134.1230 ;
      RECT 0.2600 132.9230 1704.0400 133.4770 ;
      RECT 0.0000 132.2770 1704.3000 132.9230 ;
      RECT 0.2600 131.7230 1704.0400 132.2770 ;
      RECT 0.0000 131.0770 1704.3000 131.7230 ;
      RECT 0.2600 130.5230 1704.0400 131.0770 ;
      RECT 0.0000 129.8770 1704.3000 130.5230 ;
      RECT 0.2600 129.3230 1704.0400 129.8770 ;
      RECT 0.0000 128.6770 1704.3000 129.3230 ;
      RECT 0.2600 128.1230 1704.0400 128.6770 ;
      RECT 0.0000 127.4770 1704.3000 128.1230 ;
      RECT 0.2600 126.9230 1704.0400 127.4770 ;
      RECT 0.0000 126.2770 1704.3000 126.9230 ;
      RECT 0.2600 125.7230 1704.0400 126.2770 ;
      RECT 0.0000 125.0770 1704.3000 125.7230 ;
      RECT 0.2600 124.5230 1704.0400 125.0770 ;
      RECT 0.0000 123.8770 1704.3000 124.5230 ;
      RECT 0.2600 123.3230 1704.0400 123.8770 ;
      RECT 0.0000 122.6770 1704.3000 123.3230 ;
      RECT 0.2600 122.1230 1704.0400 122.6770 ;
      RECT 0.0000 121.4770 1704.3000 122.1230 ;
      RECT 0.2600 120.9230 1704.0400 121.4770 ;
      RECT 0.0000 120.2770 1704.3000 120.9230 ;
      RECT 0.2600 119.7230 1704.0400 120.2770 ;
      RECT 0.0000 119.0770 1704.3000 119.7230 ;
      RECT 0.2600 118.5230 1704.0400 119.0770 ;
      RECT 0.0000 117.8770 1704.3000 118.5230 ;
      RECT 0.2600 117.3230 1704.0400 117.8770 ;
      RECT 0.0000 116.6770 1704.3000 117.3230 ;
      RECT 0.2600 116.1230 1704.0400 116.6770 ;
      RECT 0.0000 115.4770 1704.3000 116.1230 ;
      RECT 0.2600 114.9230 1704.0400 115.4770 ;
      RECT 0.0000 114.2770 1704.3000 114.9230 ;
      RECT 0.2600 113.7230 1704.0400 114.2770 ;
      RECT 0.0000 113.0770 1704.3000 113.7230 ;
      RECT 0.2600 112.5230 1704.0400 113.0770 ;
      RECT 0.0000 111.8770 1704.3000 112.5230 ;
      RECT 0.2600 111.3230 1704.0400 111.8770 ;
      RECT 0.0000 110.6770 1704.3000 111.3230 ;
      RECT 0.2600 110.1230 1704.0400 110.6770 ;
      RECT 0.0000 109.4770 1704.3000 110.1230 ;
      RECT 0.2600 108.9230 1704.0400 109.4770 ;
      RECT 0.0000 108.2770 1704.3000 108.9230 ;
      RECT 0.2600 107.7230 1704.0400 108.2770 ;
      RECT 0.0000 107.0770 1704.3000 107.7230 ;
      RECT 0.2600 106.5230 1704.0400 107.0770 ;
      RECT 0.0000 105.8770 1704.3000 106.5230 ;
      RECT 0.2600 105.3230 1704.0400 105.8770 ;
      RECT 0.0000 104.6770 1704.3000 105.3230 ;
      RECT 0.2600 104.1230 1704.0400 104.6770 ;
      RECT 0.0000 103.4770 1704.3000 104.1230 ;
      RECT 0.2600 102.9230 1704.0400 103.4770 ;
      RECT 0.0000 102.2770 1704.3000 102.9230 ;
      RECT 0.2600 101.7230 1704.0400 102.2770 ;
      RECT 0.0000 101.0770 1704.3000 101.7230 ;
      RECT 0.2600 100.5230 1704.0400 101.0770 ;
      RECT 0.0000 99.8770 1704.3000 100.5230 ;
      RECT 0.2600 99.3230 1704.0400 99.8770 ;
      RECT 0.0000 98.6770 1704.3000 99.3230 ;
      RECT 0.2600 98.1230 1704.0400 98.6770 ;
      RECT 0.0000 97.4770 1704.3000 98.1230 ;
      RECT 0.2600 96.9230 1704.0400 97.4770 ;
      RECT 0.0000 96.2770 1704.3000 96.9230 ;
      RECT 0.2600 95.7230 1704.0400 96.2770 ;
      RECT 0.0000 95.0770 1704.3000 95.7230 ;
      RECT 0.2600 94.5230 1704.0400 95.0770 ;
      RECT 0.0000 93.8770 1704.3000 94.5230 ;
      RECT 0.2600 93.3230 1704.0400 93.8770 ;
      RECT 0.0000 92.6770 1704.3000 93.3230 ;
      RECT 0.2600 92.1230 1704.0400 92.6770 ;
      RECT 0.0000 91.4770 1704.3000 92.1230 ;
      RECT 0.2600 90.9230 1704.0400 91.4770 ;
      RECT 0.0000 90.2770 1704.3000 90.9230 ;
      RECT 0.2600 89.7230 1704.0400 90.2770 ;
      RECT 0.0000 89.0770 1704.3000 89.7230 ;
      RECT 0.2600 88.5230 1704.0400 89.0770 ;
      RECT 0.0000 87.8770 1704.3000 88.5230 ;
      RECT 0.2600 87.3230 1704.0400 87.8770 ;
      RECT 0.0000 86.6770 1704.3000 87.3230 ;
      RECT 0.2600 86.1230 1704.0400 86.6770 ;
      RECT 0.0000 85.4770 1704.3000 86.1230 ;
      RECT 0.2600 84.9230 1704.0400 85.4770 ;
      RECT 0.0000 84.2770 1704.3000 84.9230 ;
      RECT 0.2600 83.7230 1704.0400 84.2770 ;
      RECT 0.0000 83.0770 1704.3000 83.7230 ;
      RECT 0.2600 82.5230 1704.0400 83.0770 ;
      RECT 0.0000 81.8770 1704.3000 82.5230 ;
      RECT 0.2600 81.3230 1704.0400 81.8770 ;
      RECT 0.0000 80.6770 1704.3000 81.3230 ;
      RECT 0.2600 80.1230 1704.0400 80.6770 ;
      RECT 0.0000 79.4770 1704.3000 80.1230 ;
      RECT 0.2600 78.9230 1704.0400 79.4770 ;
      RECT 0.0000 78.2770 1704.3000 78.9230 ;
      RECT 0.2600 77.7230 1704.0400 78.2770 ;
      RECT 0.0000 77.0770 1704.3000 77.7230 ;
      RECT 0.2600 76.5230 1704.0400 77.0770 ;
      RECT 0.0000 75.8770 1704.3000 76.5230 ;
      RECT 0.2600 75.3230 1704.0400 75.8770 ;
      RECT 0.0000 74.6770 1704.3000 75.3230 ;
      RECT 0.2600 74.1230 1704.0400 74.6770 ;
      RECT 0.0000 73.4770 1704.3000 74.1230 ;
      RECT 0.2600 72.9230 1704.0400 73.4770 ;
      RECT 0.0000 72.2770 1704.3000 72.9230 ;
      RECT 0.2600 71.7230 1704.0400 72.2770 ;
      RECT 0.0000 71.0770 1704.3000 71.7230 ;
      RECT 0.2600 70.5230 1704.0400 71.0770 ;
      RECT 0.0000 69.8770 1704.3000 70.5230 ;
      RECT 0.2600 69.3230 1704.0400 69.8770 ;
      RECT 0.0000 68.6770 1704.3000 69.3230 ;
      RECT 0.2600 68.1230 1704.0400 68.6770 ;
      RECT 0.0000 67.4770 1704.3000 68.1230 ;
      RECT 0.2600 66.9230 1704.0400 67.4770 ;
      RECT 0.0000 66.2770 1704.3000 66.9230 ;
      RECT 0.2600 65.7230 1704.0400 66.2770 ;
      RECT 0.0000 65.0770 1704.3000 65.7230 ;
      RECT 0.2600 64.5230 1704.0400 65.0770 ;
      RECT 0.0000 63.8770 1704.3000 64.5230 ;
      RECT 0.2600 63.3230 1704.0400 63.8770 ;
      RECT 0.0000 62.6770 1704.3000 63.3230 ;
      RECT 0.2600 62.1230 1704.0400 62.6770 ;
      RECT 0.0000 61.4770 1704.3000 62.1230 ;
      RECT 0.2600 60.9230 1704.0400 61.4770 ;
      RECT 0.0000 60.2770 1704.3000 60.9230 ;
      RECT 0.2600 59.7230 1704.0400 60.2770 ;
      RECT 0.0000 59.0770 1704.3000 59.7230 ;
      RECT 0.2600 58.5230 1704.0400 59.0770 ;
      RECT 0.0000 57.8770 1704.3000 58.5230 ;
      RECT 0.2600 57.3230 1704.0400 57.8770 ;
      RECT 0.0000 56.6770 1704.3000 57.3230 ;
      RECT 0.2600 56.1230 1704.0400 56.6770 ;
      RECT 0.0000 55.4770 1704.3000 56.1230 ;
      RECT 0.2600 54.9230 1704.0400 55.4770 ;
      RECT 0.0000 54.2770 1704.3000 54.9230 ;
      RECT 0.2600 53.7230 1704.0400 54.2770 ;
      RECT 0.0000 53.0770 1704.3000 53.7230 ;
      RECT 0.2600 52.5230 1704.0400 53.0770 ;
      RECT 0.0000 51.8770 1704.3000 52.5230 ;
      RECT 0.2600 51.3230 1704.0400 51.8770 ;
      RECT 0.0000 50.6770 1704.3000 51.3230 ;
      RECT 0.2600 50.1230 1704.0400 50.6770 ;
      RECT 0.0000 49.4770 1704.3000 50.1230 ;
      RECT 0.2600 48.9230 1704.0400 49.4770 ;
      RECT 0.0000 48.2770 1704.3000 48.9230 ;
      RECT 0.2600 47.7230 1704.0400 48.2770 ;
      RECT 0.0000 47.0770 1704.3000 47.7230 ;
      RECT 0.2600 46.5230 1704.0400 47.0770 ;
      RECT 0.0000 45.8770 1704.3000 46.5230 ;
      RECT 0.2600 45.3230 1704.0400 45.8770 ;
      RECT 0.0000 44.6770 1704.3000 45.3230 ;
      RECT 0.2600 44.1230 1704.0400 44.6770 ;
      RECT 0.0000 43.4770 1704.3000 44.1230 ;
      RECT 0.2600 42.9230 1704.0400 43.4770 ;
      RECT 0.0000 42.2770 1704.3000 42.9230 ;
      RECT 0.2600 41.7230 1704.0400 42.2770 ;
      RECT 0.0000 41.0770 1704.3000 41.7230 ;
      RECT 0.2600 40.5230 1704.0400 41.0770 ;
      RECT 0.0000 39.8770 1704.3000 40.5230 ;
      RECT 0.2600 39.3230 1704.0400 39.8770 ;
      RECT 0.0000 38.6770 1704.3000 39.3230 ;
      RECT 0.2600 38.1230 1704.0400 38.6770 ;
      RECT 0.0000 37.4770 1704.3000 38.1230 ;
      RECT 0.2600 36.9230 1704.0400 37.4770 ;
      RECT 0.0000 36.2770 1704.3000 36.9230 ;
      RECT 0.2600 35.7230 1704.0400 36.2770 ;
      RECT 0.0000 35.0770 1704.3000 35.7230 ;
      RECT 0.2600 34.5230 1704.0400 35.0770 ;
      RECT 0.0000 33.8770 1704.3000 34.5230 ;
      RECT 0.2600 33.3230 1704.0400 33.8770 ;
      RECT 0.0000 32.6770 1704.3000 33.3230 ;
      RECT 0.2600 32.1230 1704.0400 32.6770 ;
      RECT 0.0000 31.4770 1704.3000 32.1230 ;
      RECT 0.2600 30.9230 1704.0400 31.4770 ;
      RECT 0.0000 30.2770 1704.3000 30.9230 ;
      RECT 0.2600 29.7230 1704.0400 30.2770 ;
      RECT 0.0000 29.0770 1704.3000 29.7230 ;
      RECT 0.2600 28.5230 1704.0400 29.0770 ;
      RECT 0.0000 27.8770 1704.3000 28.5230 ;
      RECT 0.2600 27.3230 1704.0400 27.8770 ;
      RECT 0.0000 26.6770 1704.3000 27.3230 ;
      RECT 0.2600 26.1230 1704.0400 26.6770 ;
      RECT 0.0000 25.4770 1704.3000 26.1230 ;
      RECT 0.2600 24.9230 1704.0400 25.4770 ;
      RECT 0.0000 24.2770 1704.3000 24.9230 ;
      RECT 0.2600 23.7230 1704.0400 24.2770 ;
      RECT 0.0000 23.0770 1704.3000 23.7230 ;
      RECT 0.2600 22.5230 1704.0400 23.0770 ;
      RECT 0.0000 21.8770 1704.3000 22.5230 ;
      RECT 0.2600 21.3230 1704.0400 21.8770 ;
      RECT 0.0000 20.6770 1704.3000 21.3230 ;
      RECT 0.2600 20.1230 1704.0400 20.6770 ;
      RECT 0.0000 19.4770 1704.3000 20.1230 ;
      RECT 0.2600 18.9230 1704.0400 19.4770 ;
      RECT 0.0000 18.2770 1704.3000 18.9230 ;
      RECT 0.2600 17.7230 1704.0400 18.2770 ;
      RECT 0.0000 17.0770 1704.3000 17.7230 ;
      RECT 0.2600 16.5230 1704.0400 17.0770 ;
      RECT 0.0000 15.8770 1704.3000 16.5230 ;
      RECT 0.2600 15.3230 1704.0400 15.8770 ;
      RECT 0.0000 14.6770 1704.3000 15.3230 ;
      RECT 0.2600 14.1230 1704.0400 14.6770 ;
      RECT 0.0000 13.4770 1704.3000 14.1230 ;
      RECT 0.2600 12.9230 1704.0400 13.4770 ;
      RECT 0.0000 12.2770 1704.3000 12.9230 ;
      RECT 0.2600 11.7230 1704.0400 12.2770 ;
      RECT 0.0000 11.0770 1704.3000 11.7230 ;
      RECT 0.2600 10.5230 1704.0400 11.0770 ;
      RECT 0.0000 9.8770 1704.3000 10.5230 ;
      RECT 0.2600 9.3230 1704.0400 9.8770 ;
      RECT 0.0000 8.6770 1704.3000 9.3230 ;
      RECT 0.2600 8.1230 1704.0400 8.6770 ;
      RECT 0.0000 7.4770 1704.3000 8.1230 ;
      RECT 0.2600 6.9230 1704.0400 7.4770 ;
      RECT 0.0000 6.2770 1704.3000 6.9230 ;
      RECT 0.2600 5.7230 1704.0400 6.2770 ;
      RECT 0.0000 5.0770 1704.3000 5.7230 ;
      RECT 0.2600 4.5230 1704.0400 5.0770 ;
      RECT 0.0000 3.8770 1704.3000 4.5230 ;
      RECT 0.2600 3.3230 1704.0400 3.8770 ;
      RECT 0.0000 2.6770 1704.3000 3.3230 ;
      RECT 0.2600 2.1230 1704.0400 2.6770 ;
      RECT 0.0000 1.4770 1704.3000 2.1230 ;
      RECT 0.2600 0.9230 1704.0400 1.4770 ;
      RECT 0.0000 0.2770 1704.3000 0.9230 ;
      RECT 0.2600 0.0000 1704.0400 0.2770 ;
    LAYER M3 ;
      RECT 1703.9450 640.3700 1704.3000 640.8000 ;
      RECT 0.0000 640.3700 1701.0750 640.8000 ;
      RECT 0.0000 0.4300 1704.3000 640.3700 ;
      RECT 1703.9450 0.0000 1704.3000 0.4300 ;
      RECT 977.0450 0.0000 1703.0750 0.4300 ;
      RECT 970.6450 0.0000 973.9750 0.4300 ;
      RECT 946.6450 0.0000 949.9750 0.4300 ;
      RECT 922.6450 0.0000 925.9750 0.4300 ;
      RECT 898.6450 0.0000 901.9750 0.4300 ;
      RECT 874.3450 0.0000 877.5750 0.4300 ;
      RECT 850.0450 0.0000 853.2750 0.4300 ;
      RECT 825.7450 0.0000 828.9750 0.4300 ;
      RECT 801.4450 0.0000 804.6750 0.4300 ;
      RECT 777.1450 0.0000 780.3750 0.4300 ;
      RECT 752.7450 0.0000 756.0750 0.4300 ;
      RECT 728.4450 0.0000 731.8750 0.4300 ;
      RECT 704.1450 0.0000 707.5750 0.4300 ;
      RECT 51.9450 0.0000 703.4750 0.4300 ;
      RECT 8.7450 0.0000 51.4750 0.4300 ;
      RECT 2.9450 0.0000 8.2750 0.4300 ;
      RECT 1.6450 0.0000 2.0750 0.4300 ;
      RECT 1.0450 0.0000 1.1750 0.4300 ;
      RECT 0.0000 0.0000 0.2750 0.4300 ;
    LAYER M4 ;
      RECT 0.0000 640.4850 1704.3000 640.8000 ;
      RECT 0.0000 637.4150 1703.8700 640.4850 ;
      RECT 0.0000 430.3850 1704.3000 637.4150 ;
      RECT 0.4300 429.9150 1704.3000 430.3850 ;
      RECT 0.0000 272.8850 1704.3000 429.9150 ;
      RECT 0.4300 272.4150 1704.3000 272.8850 ;
      RECT 0.0000 208.0850 1704.3000 272.4150 ;
      RECT 0.0000 207.6150 1703.8700 208.0850 ;
      RECT 0.0000 191.2850 1704.3000 207.6150 ;
      RECT 0.0000 190.8150 1703.8700 191.2850 ;
      RECT 0.0000 163.6850 1704.3000 190.8150 ;
      RECT 0.0000 163.2150 1703.8700 163.6850 ;
      RECT 0.0000 160.7850 1704.3000 163.2150 ;
      RECT 0.0000 160.3150 1703.8700 160.7850 ;
      RECT 0.0000 160.0850 1704.3000 160.3150 ;
      RECT 0.0000 159.6150 1703.8700 160.0850 ;
      RECT 0.0000 115.3850 1704.3000 159.6150 ;
      RECT 0.4300 114.9150 1704.3000 115.3850 ;
      RECT 0.0000 3.5850 1704.3000 114.9150 ;
      RECT 0.4300 3.1150 1704.3000 3.5850 ;
      RECT 0.0000 1.6850 1704.3000 3.1150 ;
      RECT 0.4300 1.2150 1704.3000 1.6850 ;
      RECT 0.0000 1.1850 1704.3000 1.2150 ;
      RECT 0.0000 0.3150 1703.8700 1.1850 ;
      RECT 0.0000 0.0000 1704.3000 0.3150 ;
    LAYER M5 ;
      RECT 1703.9450 640.3700 1704.3000 640.8000 ;
      RECT 0.0000 640.3700 1701.0750 640.8000 ;
      RECT 0.0000 0.4300 1704.3000 640.3700 ;
      RECT 1703.9450 0.0000 1704.3000 0.4300 ;
      RECT 51.9450 0.0000 1703.2750 0.4300 ;
      RECT 0.0000 0.0000 51.4750 0.4300 ;
    LAYER M6 ;
      RECT 0.0000 640.4850 1704.3000 640.8000 ;
      RECT 0.0000 637.6150 1703.8700 640.4850 ;
      RECT 0.0000 1.1850 1704.3000 637.6150 ;
      RECT 0.0000 0.3150 1703.8700 1.1850 ;
      RECT 0.0000 0.0000 1704.3000 0.3150 ;
    LAYER B1 ;
      RECT 1703.5600 640.1500 1704.3000 640.8000 ;
      RECT 0.0000 640.1500 1700.9600 640.8000 ;
      RECT 0.0000 0.6500 1704.3000 640.1500 ;
      RECT 1556.1600 0.0000 1704.3000 0.6500 ;
      RECT 0.0000 0.0000 1555.5600 0.6500 ;
    LAYER B2 ;
      RECT 0.0000 0.0000 1704.3000 640.8000 ;
    LAYER IA ;
      RECT 1703.6920 638.4000 1704.3000 640.8000 ;
      RECT 1691.5370 638.4000 1692.6920 640.8000 ;
      RECT 1679.3820 638.4000 1680.5370 640.8000 ;
      RECT 1667.2270 638.4000 1668.3820 640.8000 ;
      RECT 1655.0720 638.4000 1656.2270 640.8000 ;
      RECT 1642.9170 638.4000 1644.0720 640.8000 ;
      RECT 1630.7620 638.4000 1631.9170 640.8000 ;
      RECT 1618.6070 638.4000 1619.7620 640.8000 ;
      RECT 1606.4520 638.4000 1607.6070 640.8000 ;
      RECT 1594.2970 638.4000 1595.4520 640.8000 ;
      RECT 1582.1420 638.4000 1583.2970 640.8000 ;
      RECT 1569.9870 638.4000 1571.1420 640.8000 ;
      RECT 1557.8320 638.4000 1558.9870 640.8000 ;
      RECT 1545.6770 638.4000 1546.8320 640.8000 ;
      RECT 1533.5220 638.4000 1534.6770 640.8000 ;
      RECT 1521.3670 638.4000 1522.5220 640.8000 ;
      RECT 1509.2120 638.4000 1510.3670 640.8000 ;
      RECT 1497.0570 638.4000 1498.2120 640.8000 ;
      RECT 1484.9020 638.4000 1486.0570 640.8000 ;
      RECT 1472.9020 638.4000 1473.9020 640.8000 ;
      RECT 1460.9020 638.4000 1461.9020 640.8000 ;
      RECT 1448.9020 638.4000 1449.9020 640.8000 ;
      RECT 1436.9020 638.4000 1437.9020 640.8000 ;
      RECT 1424.9020 638.4000 1425.9020 640.8000 ;
      RECT 1412.9020 638.4000 1413.9020 640.8000 ;
      RECT 1400.9020 638.4000 1401.9020 640.8000 ;
      RECT 1388.9020 638.4000 1389.9020 640.8000 ;
      RECT 1376.9020 638.4000 1377.9020 640.8000 ;
      RECT 1364.9020 638.4000 1365.9020 640.8000 ;
      RECT 1352.9020 638.4000 1353.9020 640.8000 ;
      RECT 1340.9020 638.4000 1341.9020 640.8000 ;
      RECT 1328.9020 638.4000 1329.9020 640.8000 ;
      RECT 1316.9020 638.4000 1317.9020 640.8000 ;
      RECT 1304.7430 638.4000 1305.9020 640.8000 ;
      RECT 1292.5880 638.4000 1293.7430 640.8000 ;
      RECT 1280.4330 638.4000 1281.5880 640.8000 ;
      RECT 1268.2780 638.4000 1269.4330 640.8000 ;
      RECT 1256.1230 638.4000 1257.2780 640.8000 ;
      RECT 1243.9680 638.4000 1245.1230 640.8000 ;
      RECT 1231.8130 638.4000 1232.9680 640.8000 ;
      RECT 1219.6580 638.4000 1220.8130 640.8000 ;
      RECT 1207.5030 638.4000 1208.6580 640.8000 ;
      RECT 1195.3480 638.4000 1196.5030 640.8000 ;
      RECT 1183.1930 638.4000 1184.3480 640.8000 ;
      RECT 1171.0380 638.4000 1172.1930 640.8000 ;
      RECT 1158.8830 638.4000 1160.0380 640.8000 ;
      RECT 1146.7280 638.4000 1147.8830 640.8000 ;
      RECT 1134.5730 638.4000 1135.7280 640.8000 ;
      RECT 1122.4180 638.4000 1123.5730 640.8000 ;
      RECT 1110.2630 638.4000 1111.4180 640.8000 ;
      RECT 1098.1080 638.4000 1099.2630 640.8000 ;
      RECT 1085.9530 638.4000 1087.1080 640.8000 ;
      RECT 1073.7980 638.4000 1074.9530 640.8000 ;
      RECT 1061.7980 638.4000 1062.7980 640.8000 ;
      RECT 1049.7980 638.4000 1050.7980 640.8000 ;
      RECT 1037.7980 638.4000 1038.7980 640.8000 ;
      RECT 1025.7980 638.4000 1026.7980 640.8000 ;
      RECT 1013.7980 638.4000 1014.7980 640.8000 ;
      RECT 1001.7980 638.4000 1002.7980 640.8000 ;
      RECT 989.7980 638.4000 990.7980 640.8000 ;
      RECT 977.7980 638.4000 978.7980 640.8000 ;
      RECT 965.7980 638.4000 966.7980 640.8000 ;
      RECT 953.7980 638.4000 954.7980 640.8000 ;
      RECT 941.7980 638.4000 942.7980 640.8000 ;
      RECT 929.7980 638.4000 930.7980 640.8000 ;
      RECT 917.7980 638.4000 918.7980 640.8000 ;
      RECT 905.7980 638.4000 906.7980 640.8000 ;
      RECT 893.6390 638.4000 894.7980 640.8000 ;
      RECT 881.4840 638.4000 882.6390 640.8000 ;
      RECT 869.3290 638.4000 870.4840 640.8000 ;
      RECT 857.1740 638.4000 858.3290 640.8000 ;
      RECT 845.0190 638.4000 846.1740 640.8000 ;
      RECT 832.8640 638.4000 834.0190 640.8000 ;
      RECT 820.7090 638.4000 821.8640 640.8000 ;
      RECT 808.5540 638.4000 809.7090 640.8000 ;
      RECT 796.3990 638.4000 797.5540 640.8000 ;
      RECT 784.2440 638.4000 785.3990 640.8000 ;
      RECT 772.0890 638.4000 773.2440 640.8000 ;
      RECT 759.9340 638.4000 761.0890 640.8000 ;
      RECT 747.7790 638.4000 748.9340 640.8000 ;
      RECT 735.6240 638.4000 736.7790 640.8000 ;
      RECT 723.4690 638.4000 724.6240 640.8000 ;
      RECT 711.3140 638.4000 712.4690 640.8000 ;
      RECT 699.1590 638.4000 700.3140 640.8000 ;
      RECT 687.0040 638.4000 688.1590 640.8000 ;
      RECT 674.8490 638.4000 676.0040 640.8000 ;
      RECT 662.6940 638.4000 663.8490 640.8000 ;
      RECT 650.6940 638.4000 651.6940 640.8000 ;
      RECT 638.6940 638.4000 639.6940 640.8000 ;
      RECT 626.6940 638.4000 627.6940 640.8000 ;
      RECT 614.6940 638.4000 615.6940 640.8000 ;
      RECT 602.6940 638.4000 603.6940 640.8000 ;
      RECT 590.6940 638.4000 591.6940 640.8000 ;
      RECT 578.6940 638.4000 579.6940 640.8000 ;
      RECT 566.6940 638.4000 567.6940 640.8000 ;
      RECT 554.6940 638.4000 555.6940 640.8000 ;
      RECT 542.6940 638.4000 543.6940 640.8000 ;
      RECT 530.6940 638.4000 531.6940 640.8000 ;
      RECT 518.6940 638.4000 519.6940 640.8000 ;
      RECT 506.6940 638.4000 507.6940 640.8000 ;
      RECT 494.6940 638.4000 495.6940 640.8000 ;
      RECT 482.5350 638.4000 483.6940 640.8000 ;
      RECT 470.3800 638.4000 471.5350 640.8000 ;
      RECT 458.2250 638.4000 459.3800 640.8000 ;
      RECT 446.0700 638.4000 447.2250 640.8000 ;
      RECT 433.9150 638.4000 435.0700 640.8000 ;
      RECT 421.7600 638.4000 422.9150 640.8000 ;
      RECT 409.6050 638.4000 410.7600 640.8000 ;
      RECT 397.4500 638.4000 398.6050 640.8000 ;
      RECT 385.2950 638.4000 386.4500 640.8000 ;
      RECT 373.1400 638.4000 374.2950 640.8000 ;
      RECT 360.9850 638.4000 362.1400 640.8000 ;
      RECT 348.8300 638.4000 349.9850 640.8000 ;
      RECT 336.6750 638.4000 337.8300 640.8000 ;
      RECT 324.5200 638.4000 325.6750 640.8000 ;
      RECT 312.3650 638.4000 313.5200 640.8000 ;
      RECT 300.2100 638.4000 301.3650 640.8000 ;
      RECT 288.0550 638.4000 289.2100 640.8000 ;
      RECT 275.9000 638.4000 277.0550 640.8000 ;
      RECT 263.7450 638.4000 264.9000 640.8000 ;
      RECT 251.5900 638.4000 252.7450 640.8000 ;
      RECT 239.5900 638.4000 240.5900 640.8000 ;
      RECT 227.5900 638.4000 228.5900 640.8000 ;
      RECT 215.5900 638.4000 216.5900 640.8000 ;
      RECT 203.5900 638.4000 204.5900 640.8000 ;
      RECT 191.5900 638.4000 192.5900 640.8000 ;
      RECT 179.5900 638.4000 180.5900 640.8000 ;
      RECT 167.5900 638.4000 168.5900 640.8000 ;
      RECT 155.5900 638.4000 156.5900 640.8000 ;
      RECT 143.5900 638.4000 144.5900 640.8000 ;
      RECT 131.5900 638.4000 132.5900 640.8000 ;
      RECT 119.5900 638.4000 120.5900 640.8000 ;
      RECT 107.5900 638.4000 108.5900 640.8000 ;
      RECT 95.5900 638.4000 96.5900 640.8000 ;
      RECT 83.5900 638.4000 84.5900 640.8000 ;
      RECT 71.4310 638.4000 72.5900 640.8000 ;
      RECT 59.2760 638.4000 60.4310 640.8000 ;
      RECT 47.1210 638.4000 48.2760 640.8000 ;
      RECT 34.9660 638.4000 36.1210 640.8000 ;
      RECT 22.8110 638.4000 23.9660 640.8000 ;
      RECT 10.6560 638.4000 11.8110 640.8000 ;
      RECT 0.0000 2.4000 1704.3000 638.4000 ;
      RECT 1703.6920 0.0000 1704.3000 2.4000 ;
      RECT 1691.5370 0.0000 1692.6920 2.4000 ;
      RECT 1679.3820 0.0000 1680.5370 2.4000 ;
      RECT 1667.2270 0.0000 1668.3820 2.4000 ;
      RECT 1655.0720 0.0000 1656.2270 2.4000 ;
      RECT 1642.9170 0.0000 1644.0720 2.4000 ;
      RECT 1630.7620 0.0000 1631.9170 2.4000 ;
      RECT 1618.6070 0.0000 1619.7620 2.4000 ;
      RECT 1606.4520 0.0000 1607.6070 2.4000 ;
      RECT 1594.2970 0.0000 1595.4520 2.4000 ;
      RECT 1582.1420 0.0000 1583.2970 2.4000 ;
      RECT 1569.9870 0.0000 1571.1420 2.4000 ;
      RECT 1557.8320 0.0000 1558.9870 2.4000 ;
      RECT 1545.6770 0.0000 1546.8320 2.4000 ;
      RECT 1533.5220 0.0000 1534.6770 2.4000 ;
      RECT 1521.3670 0.0000 1522.5220 2.4000 ;
      RECT 1509.2120 0.0000 1510.3670 2.4000 ;
      RECT 1497.0570 0.0000 1498.2120 2.4000 ;
      RECT 1484.9020 0.0000 1486.0570 2.4000 ;
      RECT 1472.9020 0.0000 1473.9020 2.4000 ;
      RECT 1460.9020 0.0000 1461.9020 2.4000 ;
      RECT 1448.9020 0.0000 1449.9020 2.4000 ;
      RECT 1436.9020 0.0000 1437.9020 2.4000 ;
      RECT 1424.9020 0.0000 1425.9020 2.4000 ;
      RECT 1412.9020 0.0000 1413.9020 2.4000 ;
      RECT 1400.9020 0.0000 1401.9020 2.4000 ;
      RECT 1388.9020 0.0000 1389.9020 2.4000 ;
      RECT 1376.9020 0.0000 1377.9020 2.4000 ;
      RECT 1364.9020 0.0000 1365.9020 2.4000 ;
      RECT 1352.9020 0.0000 1353.9020 2.4000 ;
      RECT 1340.9020 0.0000 1341.9020 2.4000 ;
      RECT 1328.9020 0.0000 1329.9020 2.4000 ;
      RECT 1316.9020 0.0000 1317.9020 2.4000 ;
      RECT 1304.7430 0.0000 1305.9020 2.4000 ;
      RECT 1292.5880 0.0000 1293.7430 2.4000 ;
      RECT 1280.4330 0.0000 1281.5880 2.4000 ;
      RECT 1268.2780 0.0000 1269.4330 2.4000 ;
      RECT 1256.1230 0.0000 1257.2780 2.4000 ;
      RECT 1243.9680 0.0000 1245.1230 2.4000 ;
      RECT 1231.8130 0.0000 1232.9680 2.4000 ;
      RECT 1219.6580 0.0000 1220.8130 2.4000 ;
      RECT 1207.5030 0.0000 1208.6580 2.4000 ;
      RECT 1195.3480 0.0000 1196.5030 2.4000 ;
      RECT 1183.1930 0.0000 1184.3480 2.4000 ;
      RECT 1171.0380 0.0000 1172.1930 2.4000 ;
      RECT 1158.8830 0.0000 1160.0380 2.4000 ;
      RECT 1146.7280 0.0000 1147.8830 2.4000 ;
      RECT 1134.5730 0.0000 1135.7280 2.4000 ;
      RECT 1122.4180 0.0000 1123.5730 2.4000 ;
      RECT 1110.2630 0.0000 1111.4180 2.4000 ;
      RECT 1098.1080 0.0000 1099.2630 2.4000 ;
      RECT 1085.9530 0.0000 1087.1080 2.4000 ;
      RECT 1073.7980 0.0000 1074.9530 2.4000 ;
      RECT 1061.7980 0.0000 1062.7980 2.4000 ;
      RECT 1049.7980 0.0000 1050.7980 2.4000 ;
      RECT 1037.7980 0.0000 1038.7980 2.4000 ;
      RECT 1025.7980 0.0000 1026.7980 2.4000 ;
      RECT 1013.7980 0.0000 1014.7980 2.4000 ;
      RECT 1001.7980 0.0000 1002.7980 2.4000 ;
      RECT 989.7980 0.0000 990.7980 2.4000 ;
      RECT 977.7980 0.0000 978.7980 2.4000 ;
      RECT 965.7980 0.0000 966.7980 2.4000 ;
      RECT 953.7980 0.0000 954.7980 2.4000 ;
      RECT 941.7980 0.0000 942.7980 2.4000 ;
      RECT 929.7980 0.0000 930.7980 2.4000 ;
      RECT 917.7980 0.0000 918.7980 2.4000 ;
      RECT 905.7980 0.0000 906.7980 2.4000 ;
      RECT 893.6390 0.0000 894.7980 2.4000 ;
      RECT 881.4840 0.0000 882.6390 2.4000 ;
      RECT 869.3290 0.0000 870.4840 2.4000 ;
      RECT 857.1740 0.0000 858.3290 2.4000 ;
      RECT 845.0190 0.0000 846.1740 2.4000 ;
      RECT 832.8640 0.0000 834.0190 2.4000 ;
      RECT 820.7090 0.0000 821.8640 2.4000 ;
      RECT 808.5540 0.0000 809.7090 2.4000 ;
      RECT 796.3990 0.0000 797.5540 2.4000 ;
      RECT 784.2440 0.0000 785.3990 2.4000 ;
      RECT 772.0890 0.0000 773.2440 2.4000 ;
      RECT 759.9340 0.0000 761.0890 2.4000 ;
      RECT 747.7790 0.0000 748.9340 2.4000 ;
      RECT 735.6240 0.0000 736.7790 2.4000 ;
      RECT 723.4690 0.0000 724.6240 2.4000 ;
      RECT 711.3140 0.0000 712.4690 2.4000 ;
      RECT 699.1590 0.0000 700.3140 2.4000 ;
      RECT 687.0040 0.0000 688.1590 2.4000 ;
      RECT 674.8490 0.0000 676.0040 2.4000 ;
      RECT 662.6940 0.0000 663.8490 2.4000 ;
      RECT 650.6940 0.0000 651.6940 2.4000 ;
      RECT 638.6940 0.0000 639.6940 2.4000 ;
      RECT 626.6940 0.0000 627.6940 2.4000 ;
      RECT 614.6940 0.0000 615.6940 2.4000 ;
      RECT 602.6940 0.0000 603.6940 2.4000 ;
      RECT 590.6940 0.0000 591.6940 2.4000 ;
      RECT 578.6940 0.0000 579.6940 2.4000 ;
      RECT 566.6940 0.0000 567.6940 2.4000 ;
      RECT 554.6940 0.0000 555.6940 2.4000 ;
      RECT 542.6940 0.0000 543.6940 2.4000 ;
      RECT 530.6940 0.0000 531.6940 2.4000 ;
      RECT 518.6940 0.0000 519.6940 2.4000 ;
      RECT 506.6940 0.0000 507.6940 2.4000 ;
      RECT 494.6940 0.0000 495.6940 2.4000 ;
      RECT 482.5350 0.0000 483.6940 2.4000 ;
      RECT 470.3800 0.0000 471.5350 2.4000 ;
      RECT 458.2250 0.0000 459.3800 2.4000 ;
      RECT 446.0700 0.0000 447.2250 2.4000 ;
      RECT 433.9150 0.0000 435.0700 2.4000 ;
      RECT 421.7600 0.0000 422.9150 2.4000 ;
      RECT 409.6050 0.0000 410.7600 2.4000 ;
      RECT 397.4500 0.0000 398.6050 2.4000 ;
      RECT 385.2950 0.0000 386.4500 2.4000 ;
      RECT 373.1400 0.0000 374.2950 2.4000 ;
      RECT 360.9850 0.0000 362.1400 2.4000 ;
      RECT 348.8300 0.0000 349.9850 2.4000 ;
      RECT 336.6750 0.0000 337.8300 2.4000 ;
      RECT 324.5200 0.0000 325.6750 2.4000 ;
      RECT 312.3650 0.0000 313.5200 2.4000 ;
      RECT 300.2100 0.0000 301.3650 2.4000 ;
      RECT 288.0550 0.0000 289.2100 2.4000 ;
      RECT 275.9000 0.0000 277.0550 2.4000 ;
      RECT 263.7450 0.0000 264.9000 2.4000 ;
      RECT 251.5900 0.0000 252.7450 2.4000 ;
      RECT 239.5900 0.0000 240.5900 2.4000 ;
      RECT 227.5900 0.0000 228.5900 2.4000 ;
      RECT 215.5900 0.0000 216.5900 2.4000 ;
      RECT 203.5900 0.0000 204.5900 2.4000 ;
      RECT 191.5900 0.0000 192.5900 2.4000 ;
      RECT 179.5900 0.0000 180.5900 2.4000 ;
      RECT 167.5900 0.0000 168.5900 2.4000 ;
      RECT 155.5900 0.0000 156.5900 2.4000 ;
      RECT 143.5900 0.0000 144.5900 2.4000 ;
      RECT 131.5900 0.0000 132.5900 2.4000 ;
      RECT 119.5900 0.0000 120.5900 2.4000 ;
      RECT 107.5900 0.0000 108.5900 2.4000 ;
      RECT 95.5900 0.0000 96.5900 2.4000 ;
      RECT 83.5900 0.0000 84.5900 2.4000 ;
      RECT 71.4310 0.0000 72.5900 2.4000 ;
      RECT 59.2760 0.0000 60.4310 2.4000 ;
      RECT 47.1210 0.0000 48.2760 2.4000 ;
      RECT 34.9660 0.0000 36.1210 2.4000 ;
      RECT 22.8110 0.0000 23.9660 2.4000 ;
      RECT 10.6560 0.0000 11.8110 2.4000 ;
    LAYER IB ;
      RECT 0.0000 638.9100 1704.3000 640.8000 ;
      RECT 2.4000 627.9100 1701.9000 638.9100 ;
      RECT 0.0000 627.0960 1704.3000 627.9100 ;
      RECT 2.4000 616.0960 1701.9000 627.0960 ;
      RECT 0.0000 615.2820 1704.3000 616.0960 ;
      RECT 2.4000 604.2820 1701.9000 615.2820 ;
      RECT 0.0000 603.4680 1704.3000 604.2820 ;
      RECT 2.4000 592.4680 1701.9000 603.4680 ;
      RECT 0.0000 591.6540 1704.3000 592.4680 ;
      RECT 2.4000 580.6540 1701.9000 591.6540 ;
      RECT 0.0000 579.8400 1704.3000 580.6540 ;
      RECT 2.4000 568.8400 1701.9000 579.8400 ;
      RECT 0.0000 567.8400 1704.3000 568.8400 ;
      RECT 2.4000 556.8400 1701.9000 567.8400 ;
      RECT 0.0000 555.8400 1704.3000 556.8400 ;
      RECT 2.4000 544.8400 1701.9000 555.8400 ;
      RECT 0.0000 543.8400 1704.3000 544.8400 ;
      RECT 2.4000 532.8400 1701.9000 543.8400 ;
      RECT 0.0000 531.8400 1704.3000 532.8400 ;
      RECT 2.4000 520.8400 1701.9000 531.8400 ;
      RECT 0.0000 519.8400 1704.3000 520.8400 ;
      RECT 2.4000 508.8400 1701.9000 519.8400 ;
      RECT 0.0000 507.8400 1704.3000 508.8400 ;
      RECT 2.4000 496.8400 1701.9000 507.8400 ;
      RECT 0.0000 496.0180 1704.3000 496.8400 ;
      RECT 2.4000 485.0180 1701.9000 496.0180 ;
      RECT 0.0000 484.2040 1704.3000 485.0180 ;
      RECT 2.4000 473.2040 1701.9000 484.2040 ;
      RECT 0.0000 472.3900 1704.3000 473.2040 ;
      RECT 2.4000 461.3900 1701.9000 472.3900 ;
      RECT 0.0000 460.5760 1704.3000 461.3900 ;
      RECT 2.4000 449.5760 1701.9000 460.5760 ;
      RECT 0.0000 448.7620 1704.3000 449.5760 ;
      RECT 2.4000 437.7620 1701.9000 448.7620 ;
      RECT 0.0000 436.9480 1704.3000 437.7620 ;
      RECT 2.4000 425.9480 1701.9000 436.9480 ;
      RECT 0.0000 425.1340 1704.3000 425.9480 ;
      RECT 2.4000 414.1340 1701.9000 425.1340 ;
      RECT 0.0000 413.3200 1704.3000 414.1340 ;
      RECT 2.4000 402.3200 1701.9000 413.3200 ;
      RECT 0.0000 401.5060 1704.3000 402.3200 ;
      RECT 2.4000 390.5060 1701.9000 401.5060 ;
      RECT 0.0000 389.6920 1704.3000 390.5060 ;
      RECT 2.4000 378.6920 1701.9000 389.6920 ;
      RECT 0.0000 377.8780 1704.3000 378.6920 ;
      RECT 2.4000 366.8780 1701.9000 377.8780 ;
      RECT 0.0000 366.0640 1704.3000 366.8780 ;
      RECT 2.4000 355.0640 1701.9000 366.0640 ;
      RECT 0.0000 354.2500 1704.3000 355.0640 ;
      RECT 2.4000 343.2500 1701.9000 354.2500 ;
      RECT 0.0000 342.4360 1704.3000 343.2500 ;
      RECT 2.4000 331.4360 1701.9000 342.4360 ;
      RECT 0.0000 330.6220 1704.3000 331.4360 ;
      RECT 2.4000 319.6220 1701.9000 330.6220 ;
      RECT 0.0000 318.8080 1704.3000 319.6220 ;
      RECT 2.4000 307.8080 1701.9000 318.8080 ;
      RECT 0.0000 306.9940 1704.3000 307.8080 ;
      RECT 2.4000 295.9940 1701.9000 306.9940 ;
      RECT 0.0000 295.1800 1704.3000 295.9940 ;
      RECT 2.4000 284.1800 1701.9000 295.1800 ;
      RECT 0.0000 283.3660 1704.3000 284.1800 ;
      RECT 2.4000 272.3660 1701.9000 283.3660 ;
      RECT 0.0000 271.5520 1704.3000 272.3660 ;
      RECT 2.4000 260.5520 1701.9000 271.5520 ;
      RECT 0.0000 259.7380 1704.3000 260.5520 ;
      RECT 2.4000 248.7380 1701.9000 259.7380 ;
      RECT 0.0000 247.9240 1704.3000 248.7380 ;
      RECT 2.4000 236.9240 1701.9000 247.9240 ;
      RECT 0.0000 236.1100 1704.3000 236.9240 ;
      RECT 2.4000 225.1100 1701.9000 236.1100 ;
      RECT 0.0000 224.2960 1704.3000 225.1100 ;
      RECT 2.4000 213.2960 1701.9000 224.2960 ;
      RECT 0.0000 212.2960 1704.3000 213.2960 ;
      RECT 2.4000 201.2960 1701.9000 212.2960 ;
      RECT 0.0000 200.2960 1704.3000 201.2960 ;
      RECT 2.4000 189.2960 1701.9000 200.2960 ;
      RECT 0.0000 188.2960 1704.3000 189.2960 ;
      RECT 2.4000 177.2960 1701.9000 188.2960 ;
      RECT 0.0000 176.2960 1704.3000 177.2960 ;
      RECT 2.4000 165.2960 1701.9000 176.2960 ;
      RECT 0.0000 164.2960 1704.3000 165.2960 ;
      RECT 2.4000 153.2960 1701.9000 164.2960 ;
      RECT 0.0000 152.2960 1704.3000 153.2960 ;
      RECT 2.4000 141.2960 1701.9000 152.2960 ;
      RECT 0.0000 140.4740 1704.3000 141.2960 ;
      RECT 2.4000 129.4740 1701.9000 140.4740 ;
      RECT 0.0000 128.6600 1704.3000 129.4740 ;
      RECT 2.4000 117.6600 1701.9000 128.6600 ;
      RECT 0.0000 116.8460 1704.3000 117.6600 ;
      RECT 2.4000 105.8460 1701.9000 116.8460 ;
      RECT 0.0000 105.0320 1704.3000 105.8460 ;
      RECT 2.4000 94.0320 1701.9000 105.0320 ;
      RECT 0.0000 93.2180 1704.3000 94.0320 ;
      RECT 2.4000 82.2180 1701.9000 93.2180 ;
      RECT 0.0000 81.4040 1704.3000 82.2180 ;
      RECT 2.4000 70.4040 1701.9000 81.4040 ;
      RECT 0.0000 69.5900 1704.3000 70.4040 ;
      RECT 2.4000 58.5900 1701.9000 69.5900 ;
      RECT 0.0000 57.7760 1704.3000 58.5900 ;
      RECT 2.4000 46.7760 1701.9000 57.7760 ;
      RECT 0.0000 45.9620 1704.3000 46.7760 ;
      RECT 2.4000 34.9620 1701.9000 45.9620 ;
      RECT 0.0000 34.1480 1704.3000 34.9620 ;
      RECT 2.4000 23.1480 1701.9000 34.1480 ;
      RECT 0.0000 22.3340 1704.3000 23.1480 ;
      RECT 2.4000 11.3340 1701.9000 22.3340 ;
      RECT 0.0000 10.5200 1704.3000 11.3340 ;
      RECT 2.4000 0.0000 1701.9000 10.5200 ;
  END
END fe

END LIBRARY
