##
## LEF for PtnCells ;
## created by Encounter v14.28-s033_1 on Thu Jan  5 13:01:49 2017
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fe
  CLASS BLOCK ;
  FOREIGN fe 0 0 ;
  ORIGIN 0.0000 0.0000 ;
  SIZE 1704.3000 BY 640.8000 ;
  SYMMETRY X Y R90 ;
  PIN i_data_i[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.9850 0.0000 717.0350 0.2200 ;
    END
  END i_data_i[575]
  PIN i_data_i[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.1850 0.0000 717.2350 0.2200 ;
    END
  END i_data_i[574]
  PIN i_data_i[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.3850 0.0000 717.4350 0.2200 ;
    END
  END i_data_i[573]
  PIN i_data_i[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.5850 0.0000 717.6350 0.2200 ;
    END
  END i_data_i[572]
  PIN i_data_i[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.7850 0.0000 717.8350 0.2200 ;
    END
  END i_data_i[571]
  PIN i_data_i[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 717.9850 0.0000 718.0350 0.2200 ;
    END
  END i_data_i[570]
  PIN i_data_i[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.3850 0.0000 718.4350 0.2200 ;
    END
  END i_data_i[569]
  PIN i_data_i[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.5850 0.0000 718.6350 0.2200 ;
    END
  END i_data_i[568]
  PIN i_data_i[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.7850 0.0000 718.8350 0.2200 ;
    END
  END i_data_i[567]
  PIN i_data_i[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.9850 0.0000 719.0350 0.2200 ;
    END
  END i_data_i[566]
  PIN i_data_i[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.1850 0.0000 719.2350 0.2200 ;
    END
  END i_data_i[565]
  PIN i_data_i[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.3850 0.0000 719.4350 0.2200 ;
    END
  END i_data_i[564]
  PIN i_data_i[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.5850 0.0000 719.6350 0.2200 ;
    END
  END i_data_i[563]
  PIN i_data_i[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.7850 0.0000 719.8350 0.2200 ;
    END
  END i_data_i[562]
  PIN i_data_i[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 719.9850 0.0000 720.0350 0.2200 ;
    END
  END i_data_i[561]
  PIN i_data_i[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.1850 0.0000 720.2350 0.2200 ;
    END
  END i_data_i[560]
  PIN i_data_i[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.5850 0.0000 720.6350 0.2200 ;
    END
  END i_data_i[559]
  PIN i_data_i[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.7850 0.0000 720.8350 0.2200 ;
    END
  END i_data_i[558]
  PIN i_data_i[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.9850 0.0000 721.0350 0.2200 ;
    END
  END i_data_i[557]
  PIN i_data_i[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.1850 0.0000 721.2350 0.2200 ;
    END
  END i_data_i[556]
  PIN i_data_i[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.3850 0.0000 721.4350 0.2200 ;
    END
  END i_data_i[555]
  PIN i_data_i[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.5850 0.0000 721.6350 0.2200 ;
    END
  END i_data_i[554]
  PIN i_data_i[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.7850 0.0000 721.8350 0.2200 ;
    END
  END i_data_i[553]
  PIN i_data_i[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 721.9850 0.0000 722.0350 0.2200 ;
    END
  END i_data_i[552]
  PIN i_data_i[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.1850 0.0000 722.2350 0.2200 ;
    END
  END i_data_i[551]
  PIN i_data_i[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.3850 0.0000 722.4350 0.2200 ;
    END
  END i_data_i[550]
  PIN i_data_i[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.7850 0.0000 722.8350 0.2200 ;
    END
  END i_data_i[549]
  PIN i_data_i[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.9850 0.0000 723.0350 0.2200 ;
    END
  END i_data_i[548]
  PIN i_data_i[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.1850 0.0000 723.2350 0.2200 ;
    END
  END i_data_i[547]
  PIN i_data_i[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.3850 0.0000 723.4350 0.2200 ;
    END
  END i_data_i[546]
  PIN i_data_i[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.5850 0.0000 723.6350 0.2200 ;
    END
  END i_data_i[545]
  PIN i_data_i[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.7850 0.0000 723.8350 0.2200 ;
    END
  END i_data_i[544]
  PIN i_data_i[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 723.9850 0.0000 724.0350 0.2200 ;
    END
  END i_data_i[543]
  PIN i_data_i[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.1850 0.0000 724.2350 0.2200 ;
    END
  END i_data_i[542]
  PIN i_data_i[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.3850 0.0000 724.4350 0.2200 ;
    END
  END i_data_i[541]
  PIN i_data_i[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.5850 0.0000 724.6350 0.2200 ;
    END
  END i_data_i[540]
  PIN i_data_i[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.9850 0.0000 725.0350 0.2200 ;
    END
  END i_data_i[539]
  PIN i_data_i[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.1850 0.0000 725.2350 0.2200 ;
    END
  END i_data_i[538]
  PIN i_data_i[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.3850 0.0000 725.4350 0.2200 ;
    END
  END i_data_i[537]
  PIN i_data_i[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.5850 0.0000 725.6350 0.2200 ;
    END
  END i_data_i[536]
  PIN i_data_i[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.7850 0.0000 725.8350 0.2200 ;
    END
  END i_data_i[535]
  PIN i_data_i[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 725.9850 0.0000 726.0350 0.2200 ;
    END
  END i_data_i[534]
  PIN i_data_i[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.1850 0.0000 726.2350 0.2200 ;
    END
  END i_data_i[533]
  PIN i_data_i[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.3850 0.0000 726.4350 0.2200 ;
    END
  END i_data_i[532]
  PIN i_data_i[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.5850 0.0000 726.6350 0.2200 ;
    END
  END i_data_i[531]
  PIN i_data_i[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.7850 0.0000 726.8350 0.2200 ;
    END
  END i_data_i[530]
  PIN i_data_i[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.1850 0.0000 727.2350 0.2200 ;
    END
  END i_data_i[529]
  PIN i_data_i[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.3850 0.0000 727.4350 0.2200 ;
    END
  END i_data_i[528]
  PIN i_data_i[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.5850 0.0000 727.6350 0.2200 ;
    END
  END i_data_i[527]
  PIN i_data_i[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.7850 0.0000 727.8350 0.2200 ;
    END
  END i_data_i[526]
  PIN i_data_i[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 727.9850 0.0000 728.0350 0.2200 ;
    END
  END i_data_i[525]
  PIN i_data_i[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 728.1850 0.0000 728.2350 0.2200 ;
    END
  END i_data_i[524]
  PIN i_data_i[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.0850 0.0000 732.1350 0.2200 ;
    END
  END i_data_i[523]
  PIN i_data_i[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.2850 0.0000 732.3350 0.2200 ;
    END
  END i_data_i[522]
  PIN i_data_i[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.4850 0.0000 732.5350 0.2200 ;
    END
  END i_data_i[521]
  PIN i_data_i[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.6850 0.0000 732.7350 0.2200 ;
    END
  END i_data_i[520]
  PIN i_data_i[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.0850 0.0000 733.1350 0.2200 ;
    END
  END i_data_i[519]
  PIN i_data_i[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.2850 0.0000 733.3350 0.2200 ;
    END
  END i_data_i[518]
  PIN i_data_i[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.4850 0.0000 733.5350 0.2200 ;
    END
  END i_data_i[517]
  PIN i_data_i[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.6850 0.0000 733.7350 0.2200 ;
    END
  END i_data_i[516]
  PIN i_data_i[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 733.8850 0.0000 733.9350 0.2200 ;
    END
  END i_data_i[515]
  PIN i_data_i[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.0850 0.0000 734.1350 0.2200 ;
    END
  END i_data_i[514]
  PIN i_data_i[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.2850 0.0000 734.3350 0.2200 ;
    END
  END i_data_i[513]
  PIN i_data_i[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.4850 0.0000 734.5350 0.2200 ;
    END
  END i_data_i[512]
  PIN i_data_i[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.6850 0.0000 734.7350 0.2200 ;
    END
  END i_data_i[511]
  PIN i_data_i[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 734.8850 0.0000 734.9350 0.2200 ;
    END
  END i_data_i[510]
  PIN i_data_i[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.2850 0.0000 735.3350 0.2200 ;
    END
  END i_data_i[509]
  PIN i_data_i[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.4850 0.0000 735.5350 0.2200 ;
    END
  END i_data_i[508]
  PIN i_data_i[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.6850 0.0000 735.7350 0.2200 ;
    END
  END i_data_i[507]
  PIN i_data_i[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.8850 0.0000 735.9350 0.2200 ;
    END
  END i_data_i[506]
  PIN i_data_i[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.0850 0.0000 736.1350 0.2200 ;
    END
  END i_data_i[505]
  PIN i_data_i[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.2850 0.0000 736.3350 0.2200 ;
    END
  END i_data_i[504]
  PIN i_data_i[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.4850 0.0000 736.5350 0.2200 ;
    END
  END i_data_i[503]
  PIN i_data_i[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.6850 0.0000 736.7350 0.2200 ;
    END
  END i_data_i[502]
  PIN i_data_i[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 736.8850 0.0000 736.9350 0.2200 ;
    END
  END i_data_i[501]
  PIN i_data_i[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.0850 0.0000 737.1350 0.2200 ;
    END
  END i_data_i[500]
  PIN i_data_i[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.6850 0.0000 737.7350 0.2200 ;
    END
  END i_data_i[499]
  PIN i_data_i[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.8850 0.0000 737.9350 0.2200 ;
    END
  END i_data_i[498]
  PIN i_data_i[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.0850 0.0000 738.1350 0.2200 ;
    END
  END i_data_i[497]
  PIN i_data_i[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.2850 0.0000 738.3350 0.2200 ;
    END
  END i_data_i[496]
  PIN i_data_i[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.4850 0.0000 738.5350 0.2200 ;
    END
  END i_data_i[495]
  PIN i_data_i[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.6850 0.0000 738.7350 0.2200 ;
    END
  END i_data_i[494]
  PIN i_data_i[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 738.8850 0.0000 738.9350 0.2200 ;
    END
  END i_data_i[493]
  PIN i_data_i[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.0850 0.0000 739.1350 0.2200 ;
    END
  END i_data_i[492]
  PIN i_data_i[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.2850 0.0000 739.3350 0.2200 ;
    END
  END i_data_i[491]
  PIN i_data_i[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.4850 0.0000 739.5350 0.2200 ;
    END
  END i_data_i[490]
  PIN i_data_i[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.8850 0.0000 739.9350 0.2200 ;
    END
  END i_data_i[489]
  PIN i_data_i[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.0850 0.0000 740.1350 0.2200 ;
    END
  END i_data_i[488]
  PIN i_data_i[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.2850 0.0000 740.3350 0.2200 ;
    END
  END i_data_i[487]
  PIN i_data_i[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.4850 0.0000 740.5350 0.2200 ;
    END
  END i_data_i[486]
  PIN i_data_i[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.6850 0.0000 740.7350 0.2200 ;
    END
  END i_data_i[485]
  PIN i_data_i[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 740.8850 0.0000 740.9350 0.2200 ;
    END
  END i_data_i[484]
  PIN i_data_i[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.0850 0.0000 741.1350 0.2200 ;
    END
  END i_data_i[483]
  PIN i_data_i[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.2850 0.0000 741.3350 0.2200 ;
    END
  END i_data_i[482]
  PIN i_data_i[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.4850 0.0000 741.5350 0.2200 ;
    END
  END i_data_i[481]
  PIN i_data_i[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.6850 0.0000 741.7350 0.2200 ;
    END
  END i_data_i[480]
  PIN i_data_i[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.0850 0.0000 742.1350 0.2200 ;
    END
  END i_data_i[479]
  PIN i_data_i[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.2850 0.0000 742.3350 0.2200 ;
    END
  END i_data_i[478]
  PIN i_data_i[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.4850 0.0000 742.5350 0.2200 ;
    END
  END i_data_i[477]
  PIN i_data_i[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.6850 0.0000 742.7350 0.2200 ;
    END
  END i_data_i[476]
  PIN i_data_i[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 742.8850 0.0000 742.9350 0.2200 ;
    END
  END i_data_i[475]
  PIN i_data_i[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.0850 0.0000 743.1350 0.2200 ;
    END
  END i_data_i[474]
  PIN i_data_i[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.2850 0.0000 743.3350 0.2200 ;
    END
  END i_data_i[473]
  PIN i_data_i[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.4850 0.0000 743.5350 0.2200 ;
    END
  END i_data_i[472]
  PIN i_data_i[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.6850 0.0000 743.7350 0.2200 ;
    END
  END i_data_i[471]
  PIN i_data_i[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 743.8850 0.0000 743.9350 0.2200 ;
    END
  END i_data_i[470]
  PIN i_data_i[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.2850 0.0000 744.3350 0.2200 ;
    END
  END i_data_i[469]
  PIN i_data_i[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.4850 0.0000 744.5350 0.2200 ;
    END
  END i_data_i[468]
  PIN i_data_i[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.6850 0.0000 744.7350 0.2200 ;
    END
  END i_data_i[467]
  PIN i_data_i[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.8850 0.0000 744.9350 0.2200 ;
    END
  END i_data_i[466]
  PIN i_data_i[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.0850 0.0000 745.1350 0.2200 ;
    END
  END i_data_i[465]
  PIN i_data_i[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.2850 0.0000 745.3350 0.2200 ;
    END
  END i_data_i[464]
  PIN i_data_i[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.4850 0.0000 745.5350 0.2200 ;
    END
  END i_data_i[463]
  PIN i_data_i[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.6850 0.0000 745.7350 0.2200 ;
    END
  END i_data_i[462]
  PIN i_data_i[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 745.8850 0.0000 745.9350 0.2200 ;
    END
  END i_data_i[461]
  PIN i_data_i[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.0850 0.0000 746.1350 0.2200 ;
    END
  END i_data_i[460]
  PIN i_data_i[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.4850 0.0000 746.5350 0.2200 ;
    END
  END i_data_i[459]
  PIN i_data_i[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.6850 0.0000 746.7350 0.2200 ;
    END
  END i_data_i[458]
  PIN i_data_i[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.8850 0.0000 746.9350 0.2200 ;
    END
  END i_data_i[457]
  PIN i_data_i[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.0850 0.0000 747.1350 0.2200 ;
    END
  END i_data_i[456]
  PIN i_data_i[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.2850 0.0000 747.3350 0.2200 ;
    END
  END i_data_i[455]
  PIN i_data_i[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.4850 0.0000 747.5350 0.2200 ;
    END
  END i_data_i[454]
  PIN i_data_i[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.6850 0.0000 747.7350 0.2200 ;
    END
  END i_data_i[453]
  PIN i_data_i[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 747.8850 0.0000 747.9350 0.2200 ;
    END
  END i_data_i[452]
  PIN i_data_i[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.0850 0.0000 748.1350 0.2200 ;
    END
  END i_data_i[451]
  PIN i_data_i[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.2850 0.0000 748.3350 0.2200 ;
    END
  END i_data_i[450]
  PIN i_data_i[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.6850 0.0000 748.7350 0.2200 ;
    END
  END i_data_i[449]
  PIN i_data_i[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.8850 0.0000 748.9350 0.2200 ;
    END
  END i_data_i[448]
  PIN i_data_i[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.0850 0.0000 749.1350 0.2200 ;
    END
  END i_data_i[447]
  PIN i_data_i[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.2850 0.0000 749.3350 0.2200 ;
    END
  END i_data_i[446]
  PIN i_data_i[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.4850 0.0000 749.5350 0.2200 ;
    END
  END i_data_i[445]
  PIN i_data_i[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.6850 0.0000 749.7350 0.2200 ;
    END
  END i_data_i[444]
  PIN i_data_i[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 749.8850 0.0000 749.9350 0.2200 ;
    END
  END i_data_i[443]
  PIN i_data_i[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.0850 0.0000 750.1350 0.2200 ;
    END
  END i_data_i[442]
  PIN i_data_i[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.2850 0.0000 750.3350 0.2200 ;
    END
  END i_data_i[441]
  PIN i_data_i[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.4850 0.0000 750.5350 0.2200 ;
    END
  END i_data_i[440]
  PIN i_data_i[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.8850 0.0000 750.9350 0.2200 ;
    END
  END i_data_i[439]
  PIN i_data_i[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.0850 0.0000 751.1350 0.2200 ;
    END
  END i_data_i[438]
  PIN i_data_i[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.2850 0.0000 751.3350 0.2200 ;
    END
  END i_data_i[437]
  PIN i_data_i[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.4850 0.0000 751.5350 0.2200 ;
    END
  END i_data_i[436]
  PIN i_data_i[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.6850 0.0000 751.7350 0.2200 ;
    END
  END i_data_i[435]
  PIN i_data_i[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 751.8850 0.0000 751.9350 0.2200 ;
    END
  END i_data_i[434]
  PIN i_data_i[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.0850 0.0000 752.1350 0.2200 ;
    END
  END i_data_i[433]
  PIN i_data_i[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.2850 0.0000 752.3350 0.2200 ;
    END
  END i_data_i[432]
  PIN i_data_i[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 752.4850 0.0000 752.5350 0.2200 ;
    END
  END i_data_i[431]
  PIN i_data_i[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.2850 0.0000 756.3350 0.2200 ;
    END
  END i_data_i[430]
  PIN i_data_i[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.6850 0.0000 756.7350 0.2200 ;
    END
  END i_data_i[429]
  PIN i_data_i[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.8850 0.0000 756.9350 0.2200 ;
    END
  END i_data_i[428]
  PIN i_data_i[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.0850 0.0000 757.1350 0.2200 ;
    END
  END i_data_i[427]
  PIN i_data_i[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.2850 0.0000 757.3350 0.2200 ;
    END
  END i_data_i[426]
  PIN i_data_i[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.4850 0.0000 757.5350 0.2200 ;
    END
  END i_data_i[425]
  PIN i_data_i[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.6850 0.0000 757.7350 0.2200 ;
    END
  END i_data_i[424]
  PIN i_data_i[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 757.8850 0.0000 757.9350 0.2200 ;
    END
  END i_data_i[423]
  PIN i_data_i[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.0850 0.0000 758.1350 0.2200 ;
    END
  END i_data_i[422]
  PIN i_data_i[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.2850 0.0000 758.3350 0.2200 ;
    END
  END i_data_i[421]
  PIN i_data_i[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.4850 0.0000 758.5350 0.2200 ;
    END
  END i_data_i[420]
  PIN i_data_i[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.8850 0.0000 758.9350 0.2200 ;
    END
  END i_data_i[419]
  PIN i_data_i[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.0850 0.0000 759.1350 0.2200 ;
    END
  END i_data_i[418]
  PIN i_data_i[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.2850 0.0000 759.3350 0.2200 ;
    END
  END i_data_i[417]
  PIN i_data_i[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.4850 0.0000 759.5350 0.2200 ;
    END
  END i_data_i[416]
  PIN i_data_i[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.6850 0.0000 759.7350 0.2200 ;
    END
  END i_data_i[415]
  PIN i_data_i[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 759.8850 0.0000 759.9350 0.2200 ;
    END
  END i_data_i[414]
  PIN i_data_i[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.0850 0.0000 760.1350 0.2200 ;
    END
  END i_data_i[413]
  PIN i_data_i[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.2850 0.0000 760.3350 0.2200 ;
    END
  END i_data_i[412]
  PIN i_data_i[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.4850 0.0000 760.5350 0.2200 ;
    END
  END i_data_i[411]
  PIN i_data_i[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.6850 0.0000 760.7350 0.2200 ;
    END
  END i_data_i[410]
  PIN i_data_i[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.0850 0.0000 761.1350 0.2200 ;
    END
  END i_data_i[409]
  PIN i_data_i[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.2850 0.0000 761.3350 0.2200 ;
    END
  END i_data_i[408]
  PIN i_data_i[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.4850 0.0000 761.5350 0.2200 ;
    END
  END i_data_i[407]
  PIN i_data_i[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.6850 0.0000 761.7350 0.2200 ;
    END
  END i_data_i[406]
  PIN i_data_i[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 761.8850 0.0000 761.9350 0.2200 ;
    END
  END i_data_i[405]
  PIN i_data_i[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.0850 0.0000 762.1350 0.2200 ;
    END
  END i_data_i[404]
  PIN i_data_i[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.2850 0.0000 762.3350 0.2200 ;
    END
  END i_data_i[403]
  PIN i_data_i[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.4850 0.0000 762.5350 0.2200 ;
    END
  END i_data_i[402]
  PIN i_data_i[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.6850 0.0000 762.7350 0.2200 ;
    END
  END i_data_i[401]
  PIN i_data_i[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 762.8850 0.0000 762.9350 0.2200 ;
    END
  END i_data_i[400]
  PIN i_data_i[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.4850 0.0000 763.5350 0.2200 ;
    END
  END i_data_i[399]
  PIN i_data_i[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.6850 0.0000 763.7350 0.2200 ;
    END
  END i_data_i[398]
  PIN i_data_i[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.8850 0.0000 763.9350 0.2200 ;
    END
  END i_data_i[397]
  PIN i_data_i[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.0850 0.0000 764.1350 0.2200 ;
    END
  END i_data_i[396]
  PIN i_data_i[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.2850 0.0000 764.3350 0.2200 ;
    END
  END i_data_i[395]
  PIN i_data_i[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.4850 0.0000 764.5350 0.2200 ;
    END
  END i_data_i[394]
  PIN i_data_i[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.6850 0.0000 764.7350 0.2200 ;
    END
  END i_data_i[393]
  PIN i_data_i[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 764.8850 0.0000 764.9350 0.2200 ;
    END
  END i_data_i[392]
  PIN i_data_i[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.0850 0.0000 765.1350 0.2200 ;
    END
  END i_data_i[391]
  PIN i_data_i[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.2850 0.0000 765.3350 0.2200 ;
    END
  END i_data_i[390]
  PIN i_data_i[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.6850 0.0000 765.7350 0.2200 ;
    END
  END i_data_i[389]
  PIN i_data_i[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.8850 0.0000 765.9350 0.2200 ;
    END
  END i_data_i[388]
  PIN i_data_i[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.0850 0.0000 766.1350 0.2200 ;
    END
  END i_data_i[387]
  PIN i_data_i[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.2850 0.0000 766.3350 0.2200 ;
    END
  END i_data_i[386]
  PIN i_data_i[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.4850 0.0000 766.5350 0.2200 ;
    END
  END i_data_i[385]
  PIN i_data_i[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.6850 0.0000 766.7350 0.2200 ;
    END
  END i_data_i[384]
  PIN i_data_i[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 766.8850 0.0000 766.9350 0.2200 ;
    END
  END i_data_i[383]
  PIN i_data_i[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.0850 0.0000 767.1350 0.2200 ;
    END
  END i_data_i[382]
  PIN i_data_i[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.2850 0.0000 767.3350 0.2200 ;
    END
  END i_data_i[381]
  PIN i_data_i[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.4850 0.0000 767.5350 0.2200 ;
    END
  END i_data_i[380]
  PIN i_data_i[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.8850 0.0000 767.9350 0.2200 ;
    END
  END i_data_i[379]
  PIN i_data_i[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.0850 0.0000 768.1350 0.2200 ;
    END
  END i_data_i[378]
  PIN i_data_i[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.2850 0.0000 768.3350 0.2200 ;
    END
  END i_data_i[377]
  PIN i_data_i[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.4850 0.0000 768.5350 0.2200 ;
    END
  END i_data_i[376]
  PIN i_data_i[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.6850 0.0000 768.7350 0.2200 ;
    END
  END i_data_i[375]
  PIN i_data_i[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 768.8850 0.0000 768.9350 0.2200 ;
    END
  END i_data_i[374]
  PIN i_data_i[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.0850 0.0000 769.1350 0.2200 ;
    END
  END i_data_i[373]
  PIN i_data_i[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.2850 0.0000 769.3350 0.2200 ;
    END
  END i_data_i[372]
  PIN i_data_i[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.4850 0.0000 769.5350 0.2200 ;
    END
  END i_data_i[371]
  PIN i_data_i[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.6850 0.0000 769.7350 0.2200 ;
    END
  END i_data_i[370]
  PIN i_data_i[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.0850 0.0000 770.1350 0.2200 ;
    END
  END i_data_i[369]
  PIN i_data_i[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.2850 0.0000 770.3350 0.2200 ;
    END
  END i_data_i[368]
  PIN i_data_i[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.4850 0.0000 770.5350 0.2200 ;
    END
  END i_data_i[367]
  PIN i_data_i[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.6850 0.0000 770.7350 0.2200 ;
    END
  END i_data_i[366]
  PIN i_data_i[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 770.8850 0.0000 770.9350 0.2200 ;
    END
  END i_data_i[365]
  PIN i_data_i[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.0850 0.0000 771.1350 0.2200 ;
    END
  END i_data_i[364]
  PIN i_data_i[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.2850 0.0000 771.3350 0.2200 ;
    END
  END i_data_i[363]
  PIN i_data_i[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.4850 0.0000 771.5350 0.2200 ;
    END
  END i_data_i[362]
  PIN i_data_i[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.6850 0.0000 771.7350 0.2200 ;
    END
  END i_data_i[361]
  PIN i_data_i[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 771.8850 0.0000 771.9350 0.2200 ;
    END
  END i_data_i[360]
  PIN i_data_i[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.2850 0.0000 772.3350 0.2200 ;
    END
  END i_data_i[359]
  PIN i_data_i[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.4850 0.0000 772.5350 0.2200 ;
    END
  END i_data_i[358]
  PIN i_data_i[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.6850 0.0000 772.7350 0.2200 ;
    END
  END i_data_i[357]
  PIN i_data_i[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.8850 0.0000 772.9350 0.2200 ;
    END
  END i_data_i[356]
  PIN i_data_i[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.0850 0.0000 773.1350 0.2200 ;
    END
  END i_data_i[355]
  PIN i_data_i[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.2850 0.0000 773.3350 0.2200 ;
    END
  END i_data_i[354]
  PIN i_data_i[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.4850 0.0000 773.5350 0.2200 ;
    END
  END i_data_i[353]
  PIN i_data_i[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.6850 0.0000 773.7350 0.2200 ;
    END
  END i_data_i[352]
  PIN i_data_i[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 773.8850 0.0000 773.9350 0.2200 ;
    END
  END i_data_i[351]
  PIN i_data_i[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.0850 0.0000 774.1350 0.2200 ;
    END
  END i_data_i[350]
  PIN i_data_i[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.4850 0.0000 774.5350 0.2200 ;
    END
  END i_data_i[349]
  PIN i_data_i[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.6850 0.0000 774.7350 0.2200 ;
    END
  END i_data_i[348]
  PIN i_data_i[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.8850 0.0000 774.9350 0.2200 ;
    END
  END i_data_i[347]
  PIN i_data_i[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.0850 0.0000 775.1350 0.2200 ;
    END
  END i_data_i[346]
  PIN i_data_i[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.2850 0.0000 775.3350 0.2200 ;
    END
  END i_data_i[345]
  PIN i_data_i[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.4850 0.0000 775.5350 0.2200 ;
    END
  END i_data_i[344]
  PIN i_data_i[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.6850 0.0000 775.7350 0.2200 ;
    END
  END i_data_i[343]
  PIN i_data_i[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 775.8850 0.0000 775.9350 0.2200 ;
    END
  END i_data_i[342]
  PIN i_data_i[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.0850 0.0000 776.1350 0.2200 ;
    END
  END i_data_i[341]
  PIN i_data_i[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.2850 0.0000 776.3350 0.2200 ;
    END
  END i_data_i[340]
  PIN i_data_i[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.6850 0.0000 776.7350 0.2200 ;
    END
  END i_data_i[339]
  PIN i_data_i[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.8850 0.0000 776.9350 0.2200 ;
    END
  END i_data_i[338]
  PIN i_data_i[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.5850 0.0000 780.6350 0.2200 ;
    END
  END i_data_i[337]
  PIN i_data_i[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.7850 0.0000 780.8350 0.2200 ;
    END
  END i_data_i[336]
  PIN i_data_i[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 780.9850 0.0000 781.0350 0.2200 ;
    END
  END i_data_i[335]
  PIN i_data_i[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.1850 0.0000 781.2350 0.2200 ;
    END
  END i_data_i[334]
  PIN i_data_i[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.3850 0.0000 781.4350 0.2200 ;
    END
  END i_data_i[333]
  PIN i_data_i[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.5850 0.0000 781.6350 0.2200 ;
    END
  END i_data_i[332]
  PIN i_data_i[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.7850 0.0000 781.8350 0.2200 ;
    END
  END i_data_i[331]
  PIN i_data_i[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 781.9850 0.0000 782.0350 0.2200 ;
    END
  END i_data_i[330]
  PIN i_data_i[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.3850 0.0000 782.4350 0.2200 ;
    END
  END i_data_i[329]
  PIN i_data_i[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.5850 0.0000 782.6350 0.2200 ;
    END
  END i_data_i[328]
  PIN i_data_i[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.7850 0.0000 782.8350 0.2200 ;
    END
  END i_data_i[327]
  PIN i_data_i[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.9850 0.0000 783.0350 0.2200 ;
    END
  END i_data_i[326]
  PIN i_data_i[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.1850 0.0000 783.2350 0.2200 ;
    END
  END i_data_i[325]
  PIN i_data_i[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.3850 0.0000 783.4350 0.2200 ;
    END
  END i_data_i[324]
  PIN i_data_i[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.5850 0.0000 783.6350 0.2200 ;
    END
  END i_data_i[323]
  PIN i_data_i[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.7850 0.0000 783.8350 0.2200 ;
    END
  END i_data_i[322]
  PIN i_data_i[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 783.9850 0.0000 784.0350 0.2200 ;
    END
  END i_data_i[321]
  PIN i_data_i[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.1850 0.0000 784.2350 0.2200 ;
    END
  END i_data_i[320]
  PIN i_data_i[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.5850 0.0000 784.6350 0.2200 ;
    END
  END i_data_i[319]
  PIN i_data_i[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.7850 0.0000 784.8350 0.2200 ;
    END
  END i_data_i[318]
  PIN i_data_i[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.9850 0.0000 785.0350 0.2200 ;
    END
  END i_data_i[317]
  PIN i_data_i[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.1850 0.0000 785.2350 0.2200 ;
    END
  END i_data_i[316]
  PIN i_data_i[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.3850 0.0000 785.4350 0.2200 ;
    END
  END i_data_i[315]
  PIN i_data_i[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.5850 0.0000 785.6350 0.2200 ;
    END
  END i_data_i[314]
  PIN i_data_i[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.7850 0.0000 785.8350 0.2200 ;
    END
  END i_data_i[313]
  PIN i_data_i[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 785.9850 0.0000 786.0350 0.2200 ;
    END
  END i_data_i[312]
  PIN i_data_i[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.1850 0.0000 786.2350 0.2200 ;
    END
  END i_data_i[311]
  PIN i_data_i[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.3850 0.0000 786.4350 0.2200 ;
    END
  END i_data_i[310]
  PIN i_data_i[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.7850 0.0000 786.8350 0.2200 ;
    END
  END i_data_i[309]
  PIN i_data_i[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.9850 0.0000 787.0350 0.2200 ;
    END
  END i_data_i[308]
  PIN i_data_i[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.1850 0.0000 787.2350 0.2200 ;
    END
  END i_data_i[307]
  PIN i_data_i[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.3850 0.0000 787.4350 0.2200 ;
    END
  END i_data_i[306]
  PIN i_data_i[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.5850 0.0000 787.6350 0.2200 ;
    END
  END i_data_i[305]
  PIN i_data_i[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.7850 0.0000 787.8350 0.2200 ;
    END
  END i_data_i[304]
  PIN i_data_i[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 787.9850 0.0000 788.0350 0.2200 ;
    END
  END i_data_i[303]
  PIN i_data_i[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.1850 0.0000 788.2350 0.2200 ;
    END
  END i_data_i[302]
  PIN i_data_i[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.3850 0.0000 788.4350 0.2200 ;
    END
  END i_data_i[301]
  PIN i_data_i[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.5850 0.0000 788.6350 0.2200 ;
    END
  END i_data_i[300]
  PIN i_data_i[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.1850 0.0000 789.2350 0.2200 ;
    END
  END i_data_i[299]
  PIN i_data_i[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.3850 0.0000 789.4350 0.2200 ;
    END
  END i_data_i[298]
  PIN i_data_i[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.5850 0.0000 789.6350 0.2200 ;
    END
  END i_data_i[297]
  PIN i_data_i[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.7850 0.0000 789.8350 0.2200 ;
    END
  END i_data_i[296]
  PIN i_data_i[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 789.9850 0.0000 790.0350 0.2200 ;
    END
  END i_data_i[295]
  PIN i_data_i[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.1850 0.0000 790.2350 0.2200 ;
    END
  END i_data_i[294]
  PIN i_data_i[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.3850 0.0000 790.4350 0.2200 ;
    END
  END i_data_i[293]
  PIN i_data_i[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.5850 0.0000 790.6350 0.2200 ;
    END
  END i_data_i[292]
  PIN i_data_i[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.7850 0.0000 790.8350 0.2200 ;
    END
  END i_data_i[291]
  PIN i_data_i[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 790.9850 0.0000 791.0350 0.2200 ;
    END
  END i_data_i[290]
  PIN i_data_i[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.3850 0.0000 791.4350 0.2200 ;
    END
  END i_data_i[289]
  PIN i_data_i[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.5850 0.0000 791.6350 0.2200 ;
    END
  END i_data_i[288]
  PIN i_data_i[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.7850 0.0000 791.8350 0.2200 ;
    END
  END i_data_i[287]
  PIN i_data_i[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.9850 0.0000 792.0350 0.2200 ;
    END
  END i_data_i[286]
  PIN i_data_i[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.1850 0.0000 792.2350 0.2200 ;
    END
  END i_data_i[285]
  PIN i_data_i[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.3850 0.0000 792.4350 0.2200 ;
    END
  END i_data_i[284]
  PIN i_data_i[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.5850 0.0000 792.6350 0.2200 ;
    END
  END i_data_i[283]
  PIN i_data_i[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.7850 0.0000 792.8350 0.2200 ;
    END
  END i_data_i[282]
  PIN i_data_i[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 792.9850 0.0000 793.0350 0.2200 ;
    END
  END i_data_i[281]
  PIN i_data_i[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.1850 0.0000 793.2350 0.2200 ;
    END
  END i_data_i[280]
  PIN i_data_i[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.5850 0.0000 793.6350 0.2200 ;
    END
  END i_data_i[279]
  PIN i_data_i[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.7850 0.0000 793.8350 0.2200 ;
    END
  END i_data_i[278]
  PIN i_data_i[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.9850 0.0000 794.0350 0.2200 ;
    END
  END i_data_i[277]
  PIN i_data_i[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.1850 0.0000 794.2350 0.2200 ;
    END
  END i_data_i[276]
  PIN i_data_i[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.3850 0.0000 794.4350 0.2200 ;
    END
  END i_data_i[275]
  PIN i_data_i[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.5850 0.0000 794.6350 0.2200 ;
    END
  END i_data_i[274]
  PIN i_data_i[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.7850 0.0000 794.8350 0.2200 ;
    END
  END i_data_i[273]
  PIN i_data_i[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 794.9850 0.0000 795.0350 0.2200 ;
    END
  END i_data_i[272]
  PIN i_data_i[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.1850 0.0000 795.2350 0.2200 ;
    END
  END i_data_i[271]
  PIN i_data_i[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.3850 0.0000 795.4350 0.2200 ;
    END
  END i_data_i[270]
  PIN i_data_i[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.7850 0.0000 795.8350 0.2200 ;
    END
  END i_data_i[269]
  PIN i_data_i[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.9850 0.0000 796.0350 0.2200 ;
    END
  END i_data_i[268]
  PIN i_data_i[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.1850 0.0000 796.2350 0.2200 ;
    END
  END i_data_i[267]
  PIN i_data_i[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.3850 0.0000 796.4350 0.2200 ;
    END
  END i_data_i[266]
  PIN i_data_i[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.5850 0.0000 796.6350 0.2200 ;
    END
  END i_data_i[265]
  PIN i_data_i[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.7850 0.0000 796.8350 0.2200 ;
    END
  END i_data_i[264]
  PIN i_data_i[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 796.9850 0.0000 797.0350 0.2200 ;
    END
  END i_data_i[263]
  PIN i_data_i[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.1850 0.0000 797.2350 0.2200 ;
    END
  END i_data_i[262]
  PIN i_data_i[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.3850 0.0000 797.4350 0.2200 ;
    END
  END i_data_i[261]
  PIN i_data_i[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.5850 0.0000 797.6350 0.2200 ;
    END
  END i_data_i[260]
  PIN i_data_i[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.9850 0.0000 798.0350 0.2200 ;
    END
  END i_data_i[259]
  PIN i_data_i[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.1850 0.0000 798.2350 0.2200 ;
    END
  END i_data_i[258]
  PIN i_data_i[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.3850 0.0000 798.4350 0.2200 ;
    END
  END i_data_i[257]
  PIN i_data_i[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.5850 0.0000 798.6350 0.2200 ;
    END
  END i_data_i[256]
  PIN i_data_i[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.7850 0.0000 798.8350 0.2200 ;
    END
  END i_data_i[255]
  PIN i_data_i[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 798.9850 0.0000 799.0350 0.2200 ;
    END
  END i_data_i[254]
  PIN i_data_i[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.1850 0.0000 799.2350 0.2200 ;
    END
  END i_data_i[253]
  PIN i_data_i[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.3850 0.0000 799.4350 0.2200 ;
    END
  END i_data_i[252]
  PIN i_data_i[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.5850 0.0000 799.6350 0.2200 ;
    END
  END i_data_i[251]
  PIN i_data_i[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.7850 0.0000 799.8350 0.2200 ;
    END
  END i_data_i[250]
  PIN i_data_i[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.1850 0.0000 800.2350 0.2200 ;
    END
  END i_data_i[249]
  PIN i_data_i[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.3850 0.0000 800.4350 0.2200 ;
    END
  END i_data_i[248]
  PIN i_data_i[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.5850 0.0000 800.6350 0.2200 ;
    END
  END i_data_i[247]
  PIN i_data_i[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.7850 0.0000 800.8350 0.2200 ;
    END
  END i_data_i[246]
  PIN i_data_i[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 800.9850 0.0000 801.0350 0.2200 ;
    END
  END i_data_i[245]
  PIN i_data_i[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 801.1850 0.0000 801.2350 0.2200 ;
    END
  END i_data_i[244]
  PIN i_data_i[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 804.8850 0.0000 804.9350 0.2200 ;
    END
  END i_data_i[243]
  PIN i_data_i[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.0850 0.0000 805.1350 0.2200 ;
    END
  END i_data_i[242]
  PIN i_data_i[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.2850 0.0000 805.3350 0.2200 ;
    END
  END i_data_i[241]
  PIN i_data_i[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.4850 0.0000 805.5350 0.2200 ;
    END
  END i_data_i[240]
  PIN i_data_i[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.8850 0.0000 805.9350 0.2200 ;
    END
  END i_data_i[239]
  PIN i_data_i[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.0850 0.0000 806.1350 0.2200 ;
    END
  END i_data_i[238]
  PIN i_data_i[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.2850 0.0000 806.3350 0.2200 ;
    END
  END i_data_i[237]
  PIN i_data_i[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.4850 0.0000 806.5350 0.2200 ;
    END
  END i_data_i[236]
  PIN i_data_i[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.6850 0.0000 806.7350 0.2200 ;
    END
  END i_data_i[235]
  PIN i_data_i[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 806.8850 0.0000 806.9350 0.2200 ;
    END
  END i_data_i[234]
  PIN i_data_i[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.0850 0.0000 807.1350 0.2200 ;
    END
  END i_data_i[233]
  PIN i_data_i[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.2850 0.0000 807.3350 0.2200 ;
    END
  END i_data_i[232]
  PIN i_data_i[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.4850 0.0000 807.5350 0.2200 ;
    END
  END i_data_i[231]
  PIN i_data_i[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.6850 0.0000 807.7350 0.2200 ;
    END
  END i_data_i[230]
  PIN i_data_i[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.0850 0.0000 808.1350 0.2200 ;
    END
  END i_data_i[229]
  PIN i_data_i[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.2850 0.0000 808.3350 0.2200 ;
    END
  END i_data_i[228]
  PIN i_data_i[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.4850 0.0000 808.5350 0.2200 ;
    END
  END i_data_i[227]
  PIN i_data_i[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.6850 0.0000 808.7350 0.2200 ;
    END
  END i_data_i[226]
  PIN i_data_i[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 808.8850 0.0000 808.9350 0.2200 ;
    END
  END i_data_i[225]
  PIN i_data_i[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.0850 0.0000 809.1350 0.2200 ;
    END
  END i_data_i[224]
  PIN i_data_i[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.2850 0.0000 809.3350 0.2200 ;
    END
  END i_data_i[223]
  PIN i_data_i[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.4850 0.0000 809.5350 0.2200 ;
    END
  END i_data_i[222]
  PIN i_data_i[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.6850 0.0000 809.7350 0.2200 ;
    END
  END i_data_i[221]
  PIN i_data_i[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 809.8850 0.0000 809.9350 0.2200 ;
    END
  END i_data_i[220]
  PIN i_data_i[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.2850 0.0000 810.3350 0.2200 ;
    END
  END i_data_i[219]
  PIN i_data_i[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.4850 0.0000 810.5350 0.2200 ;
    END
  END i_data_i[218]
  PIN i_data_i[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.6850 0.0000 810.7350 0.2200 ;
    END
  END i_data_i[217]
  PIN i_data_i[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.8850 0.0000 810.9350 0.2200 ;
    END
  END i_data_i[216]
  PIN i_data_i[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.0850 0.0000 811.1350 0.2200 ;
    END
  END i_data_i[215]
  PIN i_data_i[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.2850 0.0000 811.3350 0.2200 ;
    END
  END i_data_i[214]
  PIN i_data_i[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.4850 0.0000 811.5350 0.2200 ;
    END
  END i_data_i[213]
  PIN i_data_i[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.6850 0.0000 811.7350 0.2200 ;
    END
  END i_data_i[212]
  PIN i_data_i[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 811.8850 0.0000 811.9350 0.2200 ;
    END
  END i_data_i[211]
  PIN i_data_i[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.0850 0.0000 812.1350 0.2200 ;
    END
  END i_data_i[210]
  PIN i_data_i[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.4850 0.0000 812.5350 0.2200 ;
    END
  END i_data_i[209]
  PIN i_data_i[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.6850 0.0000 812.7350 0.2200 ;
    END
  END i_data_i[208]
  PIN i_data_i[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.8850 0.0000 812.9350 0.2200 ;
    END
  END i_data_i[207]
  PIN i_data_i[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.0850 0.0000 813.1350 0.2200 ;
    END
  END i_data_i[206]
  PIN i_data_i[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.2850 0.0000 813.3350 0.2200 ;
    END
  END i_data_i[205]
  PIN i_data_i[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.4850 0.0000 813.5350 0.2200 ;
    END
  END i_data_i[204]
  PIN i_data_i[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.6850 0.0000 813.7350 0.2200 ;
    END
  END i_data_i[203]
  PIN i_data_i[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 813.8850 0.0000 813.9350 0.2200 ;
    END
  END i_data_i[202]
  PIN i_data_i[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.0850 0.0000 814.1350 0.2200 ;
    END
  END i_data_i[201]
  PIN i_data_i[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.2850 0.0000 814.3350 0.2200 ;
    END
  END i_data_i[200]
  PIN i_data_i[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.8850 0.0000 814.9350 0.2200 ;
    END
  END i_data_i[199]
  PIN i_data_i[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.0850 0.0000 815.1350 0.2200 ;
    END
  END i_data_i[198]
  PIN i_data_i[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.2850 0.0000 815.3350 0.2200 ;
    END
  END i_data_i[197]
  PIN i_data_i[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.4850 0.0000 815.5350 0.2200 ;
    END
  END i_data_i[196]
  PIN i_data_i[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.6850 0.0000 815.7350 0.2200 ;
    END
  END i_data_i[195]
  PIN i_data_i[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 815.8850 0.0000 815.9350 0.2200 ;
    END
  END i_data_i[194]
  PIN i_data_i[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.0850 0.0000 816.1350 0.2200 ;
    END
  END i_data_i[193]
  PIN i_data_i[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.2850 0.0000 816.3350 0.2200 ;
    END
  END i_data_i[192]
  PIN i_data_i[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.4850 0.0000 816.5350 0.2200 ;
    END
  END i_data_i[191]
  PIN i_data_i[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.6850 0.0000 816.7350 0.2200 ;
    END
  END i_data_i[190]
  PIN i_data_i[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.0850 0.0000 817.1350 0.2200 ;
    END
  END i_data_i[189]
  PIN i_data_i[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.2850 0.0000 817.3350 0.2200 ;
    END
  END i_data_i[188]
  PIN i_data_i[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.4850 0.0000 817.5350 0.2200 ;
    END
  END i_data_i[187]
  PIN i_data_i[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.6850 0.0000 817.7350 0.2200 ;
    END
  END i_data_i[186]
  PIN i_data_i[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 817.8850 0.0000 817.9350 0.2200 ;
    END
  END i_data_i[185]
  PIN i_data_i[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.0850 0.0000 818.1350 0.2200 ;
    END
  END i_data_i[184]
  PIN i_data_i[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.2850 0.0000 818.3350 0.2200 ;
    END
  END i_data_i[183]
  PIN i_data_i[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.4850 0.0000 818.5350 0.2200 ;
    END
  END i_data_i[182]
  PIN i_data_i[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.6850 0.0000 818.7350 0.2200 ;
    END
  END i_data_i[181]
  PIN i_data_i[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 818.8850 0.0000 818.9350 0.2200 ;
    END
  END i_data_i[180]
  PIN i_data_i[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.2850 0.0000 819.3350 0.2200 ;
    END
  END i_data_i[179]
  PIN i_data_i[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.4850 0.0000 819.5350 0.2200 ;
    END
  END i_data_i[178]
  PIN i_data_i[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.6850 0.0000 819.7350 0.2200 ;
    END
  END i_data_i[177]
  PIN i_data_i[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.8850 0.0000 819.9350 0.2200 ;
    END
  END i_data_i[176]
  PIN i_data_i[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.0850 0.0000 820.1350 0.2200 ;
    END
  END i_data_i[175]
  PIN i_data_i[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.2850 0.0000 820.3350 0.2200 ;
    END
  END i_data_i[174]
  PIN i_data_i[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.4850 0.0000 820.5350 0.2200 ;
    END
  END i_data_i[173]
  PIN i_data_i[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.6850 0.0000 820.7350 0.2200 ;
    END
  END i_data_i[172]
  PIN i_data_i[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 820.8850 0.0000 820.9350 0.2200 ;
    END
  END i_data_i[171]
  PIN i_data_i[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.0850 0.0000 821.1350 0.2200 ;
    END
  END i_data_i[170]
  PIN i_data_i[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.4850 0.0000 821.5350 0.2200 ;
    END
  END i_data_i[169]
  PIN i_data_i[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.6850 0.0000 821.7350 0.2200 ;
    END
  END i_data_i[168]
  PIN i_data_i[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.8850 0.0000 821.9350 0.2200 ;
    END
  END i_data_i[167]
  PIN i_data_i[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.0850 0.0000 822.1350 0.2200 ;
    END
  END i_data_i[166]
  PIN i_data_i[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.2850 0.0000 822.3350 0.2200 ;
    END
  END i_data_i[165]
  PIN i_data_i[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.4850 0.0000 822.5350 0.2200 ;
    END
  END i_data_i[164]
  PIN i_data_i[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.6850 0.0000 822.7350 0.2200 ;
    END
  END i_data_i[163]
  PIN i_data_i[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 822.8850 0.0000 822.9350 0.2200 ;
    END
  END i_data_i[162]
  PIN i_data_i[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.0850 0.0000 823.1350 0.2200 ;
    END
  END i_data_i[161]
  PIN i_data_i[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.2850 0.0000 823.3350 0.2200 ;
    END
  END i_data_i[160]
  PIN i_data_i[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.6850 0.0000 823.7350 0.2200 ;
    END
  END i_data_i[159]
  PIN i_data_i[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.8850 0.0000 823.9350 0.2200 ;
    END
  END i_data_i[158]
  PIN i_data_i[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.0850 0.0000 824.1350 0.2200 ;
    END
  END i_data_i[157]
  PIN i_data_i[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.2850 0.0000 824.3350 0.2200 ;
    END
  END i_data_i[156]
  PIN i_data_i[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.4850 0.0000 824.5350 0.2200 ;
    END
  END i_data_i[155]
  PIN i_data_i[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.6850 0.0000 824.7350 0.2200 ;
    END
  END i_data_i[154]
  PIN i_data_i[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 824.8850 0.0000 824.9350 0.2200 ;
    END
  END i_data_i[153]
  PIN i_data_i[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.0850 0.0000 825.1350 0.2200 ;
    END
  END i_data_i[152]
  PIN i_data_i[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.2850 0.0000 825.3350 0.2200 ;
    END
  END i_data_i[151]
  PIN i_data_i[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 825.4850 0.0000 825.5350 0.2200 ;
    END
  END i_data_i[150]
  PIN i_data_i[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.3850 0.0000 829.4350 0.2200 ;
    END
  END i_data_i[149]
  PIN i_data_i[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.5850 0.0000 829.6350 0.2200 ;
    END
  END i_data_i[148]
  PIN i_data_i[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.7850 0.0000 829.8350 0.2200 ;
    END
  END i_data_i[147]
  PIN i_data_i[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.9850 0.0000 830.0350 0.2200 ;
    END
  END i_data_i[146]
  PIN i_data_i[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.1850 0.0000 830.2350 0.2200 ;
    END
  END i_data_i[145]
  PIN i_data_i[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.3850 0.0000 830.4350 0.2200 ;
    END
  END i_data_i[144]
  PIN i_data_i[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.5850 0.0000 830.6350 0.2200 ;
    END
  END i_data_i[143]
  PIN i_data_i[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.7850 0.0000 830.8350 0.2200 ;
    END
  END i_data_i[142]
  PIN i_data_i[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 830.9850 0.0000 831.0350 0.2200 ;
    END
  END i_data_i[141]
  PIN i_data_i[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.1850 0.0000 831.2350 0.2200 ;
    END
  END i_data_i[140]
  PIN i_data_i[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.5850 0.0000 831.6350 0.2200 ;
    END
  END i_data_i[139]
  PIN i_data_i[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.7850 0.0000 831.8350 0.2200 ;
    END
  END i_data_i[138]
  PIN i_data_i[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.9850 0.0000 832.0350 0.2200 ;
    END
  END i_data_i[137]
  PIN i_data_i[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.1850 0.0000 832.2350 0.2200 ;
    END
  END i_data_i[136]
  PIN i_data_i[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.3850 0.0000 832.4350 0.2200 ;
    END
  END i_data_i[135]
  PIN i_data_i[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.5850 0.0000 832.6350 0.2200 ;
    END
  END i_data_i[134]
  PIN i_data_i[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.7850 0.0000 832.8350 0.2200 ;
    END
  END i_data_i[133]
  PIN i_data_i[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 832.9850 0.0000 833.0350 0.2200 ;
    END
  END i_data_i[132]
  PIN i_data_i[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.1850 0.0000 833.2350 0.2200 ;
    END
  END i_data_i[131]
  PIN i_data_i[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.3850 0.0000 833.4350 0.2200 ;
    END
  END i_data_i[130]
  PIN i_data_i[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.7850 0.0000 833.8350 0.2200 ;
    END
  END i_data_i[129]
  PIN i_data_i[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.9850 0.0000 834.0350 0.2200 ;
    END
  END i_data_i[128]
  PIN i_data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.1850 0.0000 834.2350 0.2200 ;
    END
  END i_data_i[127]
  PIN i_data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.3850 0.0000 834.4350 0.2200 ;
    END
  END i_data_i[126]
  PIN i_data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.5850 0.0000 834.6350 0.2200 ;
    END
  END i_data_i[125]
  PIN i_data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.7850 0.0000 834.8350 0.2200 ;
    END
  END i_data_i[124]
  PIN i_data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 834.9850 0.0000 835.0350 0.2200 ;
    END
  END i_data_i[123]
  PIN i_data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.1850 0.0000 835.2350 0.2200 ;
    END
  END i_data_i[122]
  PIN i_data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.3850 0.0000 835.4350 0.2200 ;
    END
  END i_data_i[121]
  PIN i_data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.5850 0.0000 835.6350 0.2200 ;
    END
  END i_data_i[120]
  PIN i_data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.9850 0.0000 836.0350 0.2200 ;
    END
  END i_data_i[119]
  PIN i_data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.1850 0.0000 836.2350 0.2200 ;
    END
  END i_data_i[118]
  PIN i_data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.3850 0.0000 836.4350 0.2200 ;
    END
  END i_data_i[117]
  PIN i_data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.5850 0.0000 836.6350 0.2200 ;
    END
  END i_data_i[116]
  PIN i_data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.7850 0.0000 836.8350 0.2200 ;
    END
  END i_data_i[115]
  PIN i_data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 836.9850 0.0000 837.0350 0.2200 ;
    END
  END i_data_i[114]
  PIN i_data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.1850 0.0000 837.2350 0.2200 ;
    END
  END i_data_i[113]
  PIN i_data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.3850 0.0000 837.4350 0.2200 ;
    END
  END i_data_i[112]
  PIN i_data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.5850 0.0000 837.6350 0.2200 ;
    END
  END i_data_i[111]
  PIN i_data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.7850 0.0000 837.8350 0.2200 ;
    END
  END i_data_i[110]
  PIN i_data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.1850 0.0000 838.2350 0.2200 ;
    END
  END i_data_i[109]
  PIN i_data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.3850 0.0000 838.4350 0.2200 ;
    END
  END i_data_i[108]
  PIN i_data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.5850 0.0000 838.6350 0.2200 ;
    END
  END i_data_i[107]
  PIN i_data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.7850 0.0000 838.8350 0.2200 ;
    END
  END i_data_i[106]
  PIN i_data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 838.9850 0.0000 839.0350 0.2200 ;
    END
  END i_data_i[105]
  PIN i_data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.1850 0.0000 839.2350 0.2200 ;
    END
  END i_data_i[104]
  PIN i_data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.3850 0.0000 839.4350 0.2200 ;
    END
  END i_data_i[103]
  PIN i_data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.5850 0.0000 839.6350 0.2200 ;
    END
  END i_data_i[102]
  PIN i_data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.7850 0.0000 839.8350 0.2200 ;
    END
  END i_data_i[101]
  PIN i_data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 839.9850 0.0000 840.0350 0.2200 ;
    END
  END i_data_i[100]
  PIN i_data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 703.8850 0.0000 703.9350 0.2200 ;
    END
  END i_data_i[99]
  PIN i_data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 707.7850 0.0000 707.8350 0.2200 ;
    END
  END i_data_i[98]
  PIN i_data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 707.9850 0.0000 708.0350 0.2200 ;
    END
  END i_data_i[97]
  PIN i_data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.1850 0.0000 708.2350 0.2200 ;
    END
  END i_data_i[96]
  PIN i_data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.3850 0.0000 708.4350 0.2200 ;
    END
  END i_data_i[95]
  PIN i_data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.5850 0.0000 708.6350 0.2200 ;
    END
  END i_data_i[94]
  PIN i_data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.7850 0.0000 708.8350 0.2200 ;
    END
  END i_data_i[93]
  PIN i_data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 708.9850 0.0000 709.0350 0.2200 ;
    END
  END i_data_i[92]
  PIN i_data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.1850 0.0000 709.2350 0.2200 ;
    END
  END i_data_i[91]
  PIN i_data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.3850 0.0000 709.4350 0.2200 ;
    END
  END i_data_i[90]
  PIN i_data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.7850 0.0000 709.8350 0.2200 ;
    END
  END i_data_i[89]
  PIN i_data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.9850 0.0000 710.0350 0.2200 ;
    END
  END i_data_i[88]
  PIN i_data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.1850 0.0000 710.2350 0.2200 ;
    END
  END i_data_i[87]
  PIN i_data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.3850 0.0000 710.4350 0.2200 ;
    END
  END i_data_i[86]
  PIN i_data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.5850 0.0000 710.6350 0.2200 ;
    END
  END i_data_i[85]
  PIN i_data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.7850 0.0000 710.8350 0.2200 ;
    END
  END i_data_i[84]
  PIN i_data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 710.9850 0.0000 711.0350 0.2200 ;
    END
  END i_data_i[83]
  PIN i_data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.1850 0.0000 711.2350 0.2200 ;
    END
  END i_data_i[82]
  PIN i_data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.3850 0.0000 711.4350 0.2200 ;
    END
  END i_data_i[81]
  PIN i_data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.5850 0.0000 711.6350 0.2200 ;
    END
  END i_data_i[80]
  PIN i_data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.9850 0.0000 712.0350 0.2200 ;
    END
  END i_data_i[79]
  PIN i_data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.1850 0.0000 712.2350 0.2200 ;
    END
  END i_data_i[78]
  PIN i_data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.3850 0.0000 712.4350 0.2200 ;
    END
  END i_data_i[77]
  PIN i_data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.5850 0.0000 712.6350 0.2200 ;
    END
  END i_data_i[76]
  PIN i_data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.7850 0.0000 712.8350 0.2200 ;
    END
  END i_data_i[75]
  PIN i_data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 712.9850 0.0000 713.0350 0.2200 ;
    END
  END i_data_i[74]
  PIN i_data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.1850 0.0000 713.2350 0.2200 ;
    END
  END i_data_i[73]
  PIN i_data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.3850 0.0000 713.4350 0.2200 ;
    END
  END i_data_i[72]
  PIN i_data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.5850 0.0000 713.6350 0.2200 ;
    END
  END i_data_i[71]
  PIN i_data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.7850 0.0000 713.8350 0.2200 ;
    END
  END i_data_i[70]
  PIN i_data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.1850 0.0000 714.2350 0.2200 ;
    END
  END i_data_i[69]
  PIN i_data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.3850 0.0000 714.4350 0.2200 ;
    END
  END i_data_i[68]
  PIN i_data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.5850 0.0000 714.6350 0.2200 ;
    END
  END i_data_i[67]
  PIN i_data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.7850 0.0000 714.8350 0.2200 ;
    END
  END i_data_i[66]
  PIN i_data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 714.9850 0.0000 715.0350 0.2200 ;
    END
  END i_data_i[65]
  PIN i_data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.1850 0.0000 715.2350 0.2200 ;
    END
  END i_data_i[64]
  PIN i_data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.3850 0.0000 715.4350 0.2200 ;
    END
  END i_data_i[63]
  PIN i_data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.5850 0.0000 715.6350 0.2200 ;
    END
  END i_data_i[62]
  PIN i_data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.7850 0.0000 715.8350 0.2200 ;
    END
  END i_data_i[61]
  PIN i_data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 715.9850 0.0000 716.0350 0.2200 ;
    END
  END i_data_i[60]
  PIN i_data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.3850 0.0000 716.4350 0.2200 ;
    END
  END i_data_i[59]
  PIN i_data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.5850 0.0000 716.6350 0.2200 ;
    END
  END i_data_i[58]
  PIN i_data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.7850 0.0000 716.8350 0.2200 ;
    END
  END i_data_i[57]
  PIN i_data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 718.1850 0.0000 718.2350 0.2200 ;
    END
  END i_data_i[56]
  PIN i_data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 720.3850 0.0000 720.4350 0.2200 ;
    END
  END i_data_i[55]
  PIN i_data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 722.5850 0.0000 722.6350 0.2200 ;
    END
  END i_data_i[54]
  PIN i_data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 724.7850 0.0000 724.8350 0.2200 ;
    END
  END i_data_i[53]
  PIN i_data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 726.9850 0.0000 727.0350 0.2200 ;
    END
  END i_data_i[52]
  PIN i_data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 732.8850 0.0000 732.9350 0.2200 ;
    END
  END i_data_i[51]
  PIN i_data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 735.0850 0.0000 735.1350 0.2200 ;
    END
  END i_data_i[50]
  PIN i_data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.4850 0.0000 737.5350 0.2200 ;
    END
  END i_data_i[49]
  PIN i_data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 739.6850 0.0000 739.7350 0.2200 ;
    END
  END i_data_i[48]
  PIN i_data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 741.8850 0.0000 741.9350 0.2200 ;
    END
  END i_data_i[47]
  PIN i_data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 744.0850 0.0000 744.1350 0.2200 ;
    END
  END i_data_i[46]
  PIN i_data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 746.2850 0.0000 746.3350 0.2200 ;
    END
  END i_data_i[45]
  PIN i_data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 748.4850 0.0000 748.5350 0.2200 ;
    END
  END i_data_i[44]
  PIN i_data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 750.6850 0.0000 750.7350 0.2200 ;
    END
  END i_data_i[43]
  PIN i_data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 756.4850 0.0000 756.5350 0.2200 ;
    END
  END i_data_i[42]
  PIN i_data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 758.6850 0.0000 758.7350 0.2200 ;
    END
  END i_data_i[41]
  PIN i_data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 760.8850 0.0000 760.9350 0.2200 ;
    END
  END i_data_i[40]
  PIN i_data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.2850 0.0000 763.3350 0.2200 ;
    END
  END i_data_i[39]
  PIN i_data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 765.4850 0.0000 765.5350 0.2200 ;
    END
  END i_data_i[38]
  PIN i_data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 767.6850 0.0000 767.7350 0.2200 ;
    END
  END i_data_i[37]
  PIN i_data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 769.8850 0.0000 769.9350 0.2200 ;
    END
  END i_data_i[36]
  PIN i_data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 772.0850 0.0000 772.1350 0.2200 ;
    END
  END i_data_i[35]
  PIN i_data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 774.2850 0.0000 774.3350 0.2200 ;
    END
  END i_data_i[34]
  PIN i_data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 776.4850 0.0000 776.5350 0.2200 ;
    END
  END i_data_i[33]
  PIN i_data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 782.1850 0.0000 782.2350 0.2200 ;
    END
  END i_data_i[32]
  PIN i_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 784.3850 0.0000 784.4350 0.2200 ;
    END
  END i_data_i[31]
  PIN i_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 786.5850 0.0000 786.6350 0.2200 ;
    END
  END i_data_i[30]
  PIN i_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.9850 0.0000 789.0350 0.2200 ;
    END
  END i_data_i[29]
  PIN i_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 791.1850 0.0000 791.2350 0.2200 ;
    END
  END i_data_i[28]
  PIN i_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 793.3850 0.0000 793.4350 0.2200 ;
    END
  END i_data_i[27]
  PIN i_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 795.5850 0.0000 795.6350 0.2200 ;
    END
  END i_data_i[26]
  PIN i_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 797.7850 0.0000 797.8350 0.2200 ;
    END
  END i_data_i[25]
  PIN i_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 799.9850 0.0000 800.0350 0.2200 ;
    END
  END i_data_i[24]
  PIN i_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 805.6850 0.0000 805.7350 0.2200 ;
    END
  END i_data_i[23]
  PIN i_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 807.8850 0.0000 807.9350 0.2200 ;
    END
  END i_data_i[22]
  PIN i_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 810.0850 0.0000 810.1350 0.2200 ;
    END
  END i_data_i[21]
  PIN i_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 812.2850 0.0000 812.3350 0.2200 ;
    END
  END i_data_i[20]
  PIN i_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.6850 0.0000 814.7350 0.2200 ;
    END
  END i_data_i[19]
  PIN i_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 816.8850 0.0000 816.9350 0.2200 ;
    END
  END i_data_i[18]
  PIN i_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 819.0850 0.0000 819.1350 0.2200 ;
    END
  END i_data_i[17]
  PIN i_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 821.2850 0.0000 821.3350 0.2200 ;
    END
  END i_data_i[16]
  PIN i_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 823.4850 0.0000 823.5350 0.2200 ;
    END
  END i_data_i[15]
  PIN i_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 829.1850 0.0000 829.2350 0.2200 ;
    END
  END i_data_i[14]
  PIN i_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 831.3850 0.0000 831.4350 0.2200 ;
    END
  END i_data_i[13]
  PIN i_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 833.5850 0.0000 833.6350 0.2200 ;
    END
  END i_data_i[12]
  PIN i_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 835.7850 0.0000 835.8350 0.2200 ;
    END
  END i_data_i[11]
  PIN i_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 837.9850 0.0000 838.0350 0.2200 ;
    END
  END i_data_i[10]
  PIN i_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 703.6850 0.0000 703.7350 0.2200 ;
    END
  END i_data_i[9]
  PIN i_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 709.5850 0.0000 709.6350 0.2200 ;
    END
  END i_data_i[8]
  PIN i_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 711.7850 0.0000 711.8350 0.2200 ;
    END
  END i_data_i[7]
  PIN i_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 713.9850 0.0000 714.0350 0.2200 ;
    END
  END i_data_i[6]
  PIN i_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 716.1850 0.0000 716.2350 0.2200 ;
    END
  END i_data_i[5]
  PIN i_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 737.2850 0.0000 737.3350 0.2200 ;
    END
  END i_data_i[4]
  PIN i_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 763.0850 0.0000 763.1350 0.2200 ;
    END
  END i_data_i[3]
  PIN i_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 788.7850 0.0000 788.8350 0.2200 ;
    END
  END i_data_i[2]
  PIN i_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 814.4850 0.0000 814.5350 0.2200 ;
    END
  END i_data_i[1]
  PIN i_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.1850 0.0000 840.2350 0.2200 ;
    END
  END i_data_i[0]
  PIN i_data_q[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.5850 0.0000 963.6350 0.2200 ;
    END
  END i_data_q[575]
  PIN i_data_q[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.3850 0.0000 963.4350 0.2200 ;
    END
  END i_data_q[574]
  PIN i_data_q[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.1850 0.0000 963.2350 0.2200 ;
    END
  END i_data_q[573]
  PIN i_data_q[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.9850 0.0000 963.0350 0.2200 ;
    END
  END i_data_q[572]
  PIN i_data_q[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.7850 0.0000 962.8350 0.2200 ;
    END
  END i_data_q[571]
  PIN i_data_q[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.5850 0.0000 962.6350 0.2200 ;
    END
  END i_data_q[570]
  PIN i_data_q[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.1850 0.0000 962.2350 0.2200 ;
    END
  END i_data_q[569]
  PIN i_data_q[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.9850 0.0000 962.0350 0.2200 ;
    END
  END i_data_q[568]
  PIN i_data_q[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.7850 0.0000 961.8350 0.2200 ;
    END
  END i_data_q[567]
  PIN i_data_q[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.5850 0.0000 961.6350 0.2200 ;
    END
  END i_data_q[566]
  PIN i_data_q[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.3850 0.0000 961.4350 0.2200 ;
    END
  END i_data_q[565]
  PIN i_data_q[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 961.1850 0.0000 961.2350 0.2200 ;
    END
  END i_data_q[564]
  PIN i_data_q[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.9850 0.0000 961.0350 0.2200 ;
    END
  END i_data_q[563]
  PIN i_data_q[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.7850 0.0000 960.8350 0.2200 ;
    END
  END i_data_q[562]
  PIN i_data_q[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.5850 0.0000 960.6350 0.2200 ;
    END
  END i_data_q[561]
  PIN i_data_q[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.3850 0.0000 960.4350 0.2200 ;
    END
  END i_data_q[560]
  PIN i_data_q[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.9850 0.0000 960.0350 0.2200 ;
    END
  END i_data_q[559]
  PIN i_data_q[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.7850 0.0000 959.8350 0.2200 ;
    END
  END i_data_q[558]
  PIN i_data_q[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.5850 0.0000 959.6350 0.2200 ;
    END
  END i_data_q[557]
  PIN i_data_q[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.3850 0.0000 959.4350 0.2200 ;
    END
  END i_data_q[556]
  PIN i_data_q[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 959.1850 0.0000 959.2350 0.2200 ;
    END
  END i_data_q[555]
  PIN i_data_q[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.9850 0.0000 959.0350 0.2200 ;
    END
  END i_data_q[554]
  PIN i_data_q[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.7850 0.0000 958.8350 0.2200 ;
    END
  END i_data_q[553]
  PIN i_data_q[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.5850 0.0000 958.6350 0.2200 ;
    END
  END i_data_q[552]
  PIN i_data_q[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.3850 0.0000 958.4350 0.2200 ;
    END
  END i_data_q[551]
  PIN i_data_q[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 958.1850 0.0000 958.2350 0.2200 ;
    END
  END i_data_q[550]
  PIN i_data_q[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.7850 0.0000 957.8350 0.2200 ;
    END
  END i_data_q[549]
  PIN i_data_q[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.5850 0.0000 957.6350 0.2200 ;
    END
  END i_data_q[548]
  PIN i_data_q[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.3850 0.0000 957.4350 0.2200 ;
    END
  END i_data_q[547]
  PIN i_data_q[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.1850 0.0000 957.2350 0.2200 ;
    END
  END i_data_q[546]
  PIN i_data_q[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.9850 0.0000 957.0350 0.2200 ;
    END
  END i_data_q[545]
  PIN i_data_q[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.7850 0.0000 956.8350 0.2200 ;
    END
  END i_data_q[544]
  PIN i_data_q[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.5850 0.0000 956.6350 0.2200 ;
    END
  END i_data_q[543]
  PIN i_data_q[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.3850 0.0000 956.4350 0.2200 ;
    END
  END i_data_q[542]
  PIN i_data_q[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 956.1850 0.0000 956.2350 0.2200 ;
    END
  END i_data_q[541]
  PIN i_data_q[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.9850 0.0000 956.0350 0.2200 ;
    END
  END i_data_q[540]
  PIN i_data_q[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.5850 0.0000 955.6350 0.2200 ;
    END
  END i_data_q[539]
  PIN i_data_q[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.3850 0.0000 955.4350 0.2200 ;
    END
  END i_data_q[538]
  PIN i_data_q[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.1850 0.0000 955.2350 0.2200 ;
    END
  END i_data_q[537]
  PIN i_data_q[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.9850 0.0000 955.0350 0.2200 ;
    END
  END i_data_q[536]
  PIN i_data_q[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.7850 0.0000 954.8350 0.2200 ;
    END
  END i_data_q[535]
  PIN i_data_q[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.5850 0.0000 954.6350 0.2200 ;
    END
  END i_data_q[534]
  PIN i_data_q[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.3850 0.0000 954.4350 0.2200 ;
    END
  END i_data_q[533]
  PIN i_data_q[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 954.1850 0.0000 954.2350 0.2200 ;
    END
  END i_data_q[532]
  PIN i_data_q[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.9850 0.0000 954.0350 0.2200 ;
    END
  END i_data_q[531]
  PIN i_data_q[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.7850 0.0000 953.8350 0.2200 ;
    END
  END i_data_q[530]
  PIN i_data_q[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.3850 0.0000 953.4350 0.2200 ;
    END
  END i_data_q[529]
  PIN i_data_q[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.1850 0.0000 953.2350 0.2200 ;
    END
  END i_data_q[528]
  PIN i_data_q[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.9850 0.0000 953.0350 0.2200 ;
    END
  END i_data_q[527]
  PIN i_data_q[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.7850 0.0000 952.8350 0.2200 ;
    END
  END i_data_q[526]
  PIN i_data_q[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.5850 0.0000 952.6350 0.2200 ;
    END
  END i_data_q[525]
  PIN i_data_q[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.3850 0.0000 952.4350 0.2200 ;
    END
  END i_data_q[524]
  PIN i_data_q[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 952.1850 0.0000 952.2350 0.2200 ;
    END
  END i_data_q[523]
  PIN i_data_q[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.9850 0.0000 952.0350 0.2200 ;
    END
  END i_data_q[522]
  PIN i_data_q[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.7850 0.0000 951.8350 0.2200 ;
    END
  END i_data_q[521]
  PIN i_data_q[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.5850 0.0000 951.6350 0.2200 ;
    END
  END i_data_q[520]
  PIN i_data_q[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.1850 0.0000 951.2350 0.2200 ;
    END
  END i_data_q[519]
  PIN i_data_q[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.9850 0.0000 951.0350 0.2200 ;
    END
  END i_data_q[518]
  PIN i_data_q[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.7850 0.0000 950.8350 0.2200 ;
    END
  END i_data_q[517]
  PIN i_data_q[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.5850 0.0000 950.6350 0.2200 ;
    END
  END i_data_q[516]
  PIN i_data_q[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.3850 0.0000 950.4350 0.2200 ;
    END
  END i_data_q[515]
  PIN i_data_q[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 950.1850 0.0000 950.2350 0.2200 ;
    END
  END i_data_q[514]
  PIN i_data_q[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 946.3850 0.0000 946.4350 0.2200 ;
    END
  END i_data_q[513]
  PIN i_data_q[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 946.1850 0.0000 946.2350 0.2200 ;
    END
  END i_data_q[512]
  PIN i_data_q[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.9850 0.0000 946.0350 0.2200 ;
    END
  END i_data_q[511]
  PIN i_data_q[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.7850 0.0000 945.8350 0.2200 ;
    END
  END i_data_q[510]
  PIN i_data_q[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.3850 0.0000 945.4350 0.2200 ;
    END
  END i_data_q[509]
  PIN i_data_q[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.1850 0.0000 945.2350 0.2200 ;
    END
  END i_data_q[508]
  PIN i_data_q[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.9850 0.0000 945.0350 0.2200 ;
    END
  END i_data_q[507]
  PIN i_data_q[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.7850 0.0000 944.8350 0.2200 ;
    END
  END i_data_q[506]
  PIN i_data_q[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.5850 0.0000 944.6350 0.2200 ;
    END
  END i_data_q[505]
  PIN i_data_q[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.3850 0.0000 944.4350 0.2200 ;
    END
  END i_data_q[504]
  PIN i_data_q[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 944.1850 0.0000 944.2350 0.2200 ;
    END
  END i_data_q[503]
  PIN i_data_q[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.9850 0.0000 944.0350 0.2200 ;
    END
  END i_data_q[502]
  PIN i_data_q[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.7850 0.0000 943.8350 0.2200 ;
    END
  END i_data_q[501]
  PIN i_data_q[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.5850 0.0000 943.6350 0.2200 ;
    END
  END i_data_q[500]
  PIN i_data_q[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.9850 0.0000 943.0350 0.2200 ;
    END
  END i_data_q[499]
  PIN i_data_q[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.7850 0.0000 942.8350 0.2200 ;
    END
  END i_data_q[498]
  PIN i_data_q[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.5850 0.0000 942.6350 0.2200 ;
    END
  END i_data_q[497]
  PIN i_data_q[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.3850 0.0000 942.4350 0.2200 ;
    END
  END i_data_q[496]
  PIN i_data_q[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 942.1850 0.0000 942.2350 0.2200 ;
    END
  END i_data_q[495]
  PIN i_data_q[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.9850 0.0000 942.0350 0.2200 ;
    END
  END i_data_q[494]
  PIN i_data_q[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.7850 0.0000 941.8350 0.2200 ;
    END
  END i_data_q[493]
  PIN i_data_q[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.5850 0.0000 941.6350 0.2200 ;
    END
  END i_data_q[492]
  PIN i_data_q[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.3850 0.0000 941.4350 0.2200 ;
    END
  END i_data_q[491]
  PIN i_data_q[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 941.1850 0.0000 941.2350 0.2200 ;
    END
  END i_data_q[490]
  PIN i_data_q[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.7850 0.0000 940.8350 0.2200 ;
    END
  END i_data_q[489]
  PIN i_data_q[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.5850 0.0000 940.6350 0.2200 ;
    END
  END i_data_q[488]
  PIN i_data_q[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.3850 0.0000 940.4350 0.2200 ;
    END
  END i_data_q[487]
  PIN i_data_q[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.1850 0.0000 940.2350 0.2200 ;
    END
  END i_data_q[486]
  PIN i_data_q[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.9850 0.0000 940.0350 0.2200 ;
    END
  END i_data_q[485]
  PIN i_data_q[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.7850 0.0000 939.8350 0.2200 ;
    END
  END i_data_q[484]
  PIN i_data_q[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.5850 0.0000 939.6350 0.2200 ;
    END
  END i_data_q[483]
  PIN i_data_q[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.3850 0.0000 939.4350 0.2200 ;
    END
  END i_data_q[482]
  PIN i_data_q[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 939.1850 0.0000 939.2350 0.2200 ;
    END
  END i_data_q[481]
  PIN i_data_q[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.9850 0.0000 939.0350 0.2200 ;
    END
  END i_data_q[480]
  PIN i_data_q[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.5850 0.0000 938.6350 0.2200 ;
    END
  END i_data_q[479]
  PIN i_data_q[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.3850 0.0000 938.4350 0.2200 ;
    END
  END i_data_q[478]
  PIN i_data_q[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.1850 0.0000 938.2350 0.2200 ;
    END
  END i_data_q[477]
  PIN i_data_q[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.9850 0.0000 938.0350 0.2200 ;
    END
  END i_data_q[476]
  PIN i_data_q[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.7850 0.0000 937.8350 0.2200 ;
    END
  END i_data_q[475]
  PIN i_data_q[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.5850 0.0000 937.6350 0.2200 ;
    END
  END i_data_q[474]
  PIN i_data_q[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.3850 0.0000 937.4350 0.2200 ;
    END
  END i_data_q[473]
  PIN i_data_q[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 937.1850 0.0000 937.2350 0.2200 ;
    END
  END i_data_q[472]
  PIN i_data_q[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.9850 0.0000 937.0350 0.2200 ;
    END
  END i_data_q[471]
  PIN i_data_q[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.7850 0.0000 936.8350 0.2200 ;
    END
  END i_data_q[470]
  PIN i_data_q[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.3850 0.0000 936.4350 0.2200 ;
    END
  END i_data_q[469]
  PIN i_data_q[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.1850 0.0000 936.2350 0.2200 ;
    END
  END i_data_q[468]
  PIN i_data_q[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.9850 0.0000 936.0350 0.2200 ;
    END
  END i_data_q[467]
  PIN i_data_q[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.7850 0.0000 935.8350 0.2200 ;
    END
  END i_data_q[466]
  PIN i_data_q[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.5850 0.0000 935.6350 0.2200 ;
    END
  END i_data_q[465]
  PIN i_data_q[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.3850 0.0000 935.4350 0.2200 ;
    END
  END i_data_q[464]
  PIN i_data_q[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 935.1850 0.0000 935.2350 0.2200 ;
    END
  END i_data_q[463]
  PIN i_data_q[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.9850 0.0000 935.0350 0.2200 ;
    END
  END i_data_q[462]
  PIN i_data_q[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.7850 0.0000 934.8350 0.2200 ;
    END
  END i_data_q[461]
  PIN i_data_q[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.5850 0.0000 934.6350 0.2200 ;
    END
  END i_data_q[460]
  PIN i_data_q[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.1850 0.0000 934.2350 0.2200 ;
    END
  END i_data_q[459]
  PIN i_data_q[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.9850 0.0000 934.0350 0.2200 ;
    END
  END i_data_q[458]
  PIN i_data_q[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.7850 0.0000 933.8350 0.2200 ;
    END
  END i_data_q[457]
  PIN i_data_q[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.5850 0.0000 933.6350 0.2200 ;
    END
  END i_data_q[456]
  PIN i_data_q[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.3850 0.0000 933.4350 0.2200 ;
    END
  END i_data_q[455]
  PIN i_data_q[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 933.1850 0.0000 933.2350 0.2200 ;
    END
  END i_data_q[454]
  PIN i_data_q[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.9850 0.0000 933.0350 0.2200 ;
    END
  END i_data_q[453]
  PIN i_data_q[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.7850 0.0000 932.8350 0.2200 ;
    END
  END i_data_q[452]
  PIN i_data_q[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.5850 0.0000 932.6350 0.2200 ;
    END
  END i_data_q[451]
  PIN i_data_q[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.3850 0.0000 932.4350 0.2200 ;
    END
  END i_data_q[450]
  PIN i_data_q[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.9850 0.0000 932.0350 0.2200 ;
    END
  END i_data_q[449]
  PIN i_data_q[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.7850 0.0000 931.8350 0.2200 ;
    END
  END i_data_q[448]
  PIN i_data_q[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.5850 0.0000 931.6350 0.2200 ;
    END
  END i_data_q[447]
  PIN i_data_q[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.3850 0.0000 931.4350 0.2200 ;
    END
  END i_data_q[446]
  PIN i_data_q[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 931.1850 0.0000 931.2350 0.2200 ;
    END
  END i_data_q[445]
  PIN i_data_q[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.9850 0.0000 931.0350 0.2200 ;
    END
  END i_data_q[444]
  PIN i_data_q[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.7850 0.0000 930.8350 0.2200 ;
    END
  END i_data_q[443]
  PIN i_data_q[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.5850 0.0000 930.6350 0.2200 ;
    END
  END i_data_q[442]
  PIN i_data_q[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.3850 0.0000 930.4350 0.2200 ;
    END
  END i_data_q[441]
  PIN i_data_q[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 930.1850 0.0000 930.2350 0.2200 ;
    END
  END i_data_q[440]
  PIN i_data_q[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.7850 0.0000 929.8350 0.2200 ;
    END
  END i_data_q[439]
  PIN i_data_q[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.5850 0.0000 929.6350 0.2200 ;
    END
  END i_data_q[438]
  PIN i_data_q[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.3850 0.0000 929.4350 0.2200 ;
    END
  END i_data_q[437]
  PIN i_data_q[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.1850 0.0000 929.2350 0.2200 ;
    END
  END i_data_q[436]
  PIN i_data_q[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.9850 0.0000 929.0350 0.2200 ;
    END
  END i_data_q[435]
  PIN i_data_q[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.7850 0.0000 928.8350 0.2200 ;
    END
  END i_data_q[434]
  PIN i_data_q[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.5850 0.0000 928.6350 0.2200 ;
    END
  END i_data_q[433]
  PIN i_data_q[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.3850 0.0000 928.4350 0.2200 ;
    END
  END i_data_q[432]
  PIN i_data_q[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 928.1850 0.0000 928.2350 0.2200 ;
    END
  END i_data_q[431]
  PIN i_data_q[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.9850 0.0000 928.0350 0.2200 ;
    END
  END i_data_q[430]
  PIN i_data_q[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.5850 0.0000 927.6350 0.2200 ;
    END
  END i_data_q[429]
  PIN i_data_q[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.3850 0.0000 927.4350 0.2200 ;
    END
  END i_data_q[428]
  PIN i_data_q[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.1850 0.0000 927.2350 0.2200 ;
    END
  END i_data_q[427]
  PIN i_data_q[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.9850 0.0000 927.0350 0.2200 ;
    END
  END i_data_q[426]
  PIN i_data_q[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.7850 0.0000 926.8350 0.2200 ;
    END
  END i_data_q[425]
  PIN i_data_q[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.5850 0.0000 926.6350 0.2200 ;
    END
  END i_data_q[424]
  PIN i_data_q[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.3850 0.0000 926.4350 0.2200 ;
    END
  END i_data_q[423]
  PIN i_data_q[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 926.1850 0.0000 926.2350 0.2200 ;
    END
  END i_data_q[422]
  PIN i_data_q[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 922.3850 0.0000 922.4350 0.2200 ;
    END
  END i_data_q[421]
  PIN i_data_q[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 922.1850 0.0000 922.2350 0.2200 ;
    END
  END i_data_q[420]
  PIN i_data_q[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.7850 0.0000 921.8350 0.2200 ;
    END
  END i_data_q[419]
  PIN i_data_q[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.5850 0.0000 921.6350 0.2200 ;
    END
  END i_data_q[418]
  PIN i_data_q[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.3850 0.0000 921.4350 0.2200 ;
    END
  END i_data_q[417]
  PIN i_data_q[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.1850 0.0000 921.2350 0.2200 ;
    END
  END i_data_q[416]
  PIN i_data_q[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.9850 0.0000 921.0350 0.2200 ;
    END
  END i_data_q[415]
  PIN i_data_q[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.7850 0.0000 920.8350 0.2200 ;
    END
  END i_data_q[414]
  PIN i_data_q[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.5850 0.0000 920.6350 0.2200 ;
    END
  END i_data_q[413]
  PIN i_data_q[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.3850 0.0000 920.4350 0.2200 ;
    END
  END i_data_q[412]
  PIN i_data_q[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 920.1850 0.0000 920.2350 0.2200 ;
    END
  END i_data_q[411]
  PIN i_data_q[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.9850 0.0000 920.0350 0.2200 ;
    END
  END i_data_q[410]
  PIN i_data_q[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.5850 0.0000 919.6350 0.2200 ;
    END
  END i_data_q[409]
  PIN i_data_q[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.3850 0.0000 919.4350 0.2200 ;
    END
  END i_data_q[408]
  PIN i_data_q[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.1850 0.0000 919.2350 0.2200 ;
    END
  END i_data_q[407]
  PIN i_data_q[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.9850 0.0000 919.0350 0.2200 ;
    END
  END i_data_q[406]
  PIN i_data_q[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.7850 0.0000 918.8350 0.2200 ;
    END
  END i_data_q[405]
  PIN i_data_q[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.5850 0.0000 918.6350 0.2200 ;
    END
  END i_data_q[404]
  PIN i_data_q[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.3850 0.0000 918.4350 0.2200 ;
    END
  END i_data_q[403]
  PIN i_data_q[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 918.1850 0.0000 918.2350 0.2200 ;
    END
  END i_data_q[402]
  PIN i_data_q[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.9850 0.0000 918.0350 0.2200 ;
    END
  END i_data_q[401]
  PIN i_data_q[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.7850 0.0000 917.8350 0.2200 ;
    END
  END i_data_q[400]
  PIN i_data_q[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.1850 0.0000 917.2350 0.2200 ;
    END
  END i_data_q[399]
  PIN i_data_q[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.9850 0.0000 917.0350 0.2200 ;
    END
  END i_data_q[398]
  PIN i_data_q[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.7850 0.0000 916.8350 0.2200 ;
    END
  END i_data_q[397]
  PIN i_data_q[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.5850 0.0000 916.6350 0.2200 ;
    END
  END i_data_q[396]
  PIN i_data_q[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.3850 0.0000 916.4350 0.2200 ;
    END
  END i_data_q[395]
  PIN i_data_q[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 916.1850 0.0000 916.2350 0.2200 ;
    END
  END i_data_q[394]
  PIN i_data_q[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.9850 0.0000 916.0350 0.2200 ;
    END
  END i_data_q[393]
  PIN i_data_q[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.7850 0.0000 915.8350 0.2200 ;
    END
  END i_data_q[392]
  PIN i_data_q[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.5850 0.0000 915.6350 0.2200 ;
    END
  END i_data_q[391]
  PIN i_data_q[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.3850 0.0000 915.4350 0.2200 ;
    END
  END i_data_q[390]
  PIN i_data_q[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.9850 0.0000 915.0350 0.2200 ;
    END
  END i_data_q[389]
  PIN i_data_q[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.7850 0.0000 914.8350 0.2200 ;
    END
  END i_data_q[388]
  PIN i_data_q[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.5850 0.0000 914.6350 0.2200 ;
    END
  END i_data_q[387]
  PIN i_data_q[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.3850 0.0000 914.4350 0.2200 ;
    END
  END i_data_q[386]
  PIN i_data_q[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 914.1850 0.0000 914.2350 0.2200 ;
    END
  END i_data_q[385]
  PIN i_data_q[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.9850 0.0000 914.0350 0.2200 ;
    END
  END i_data_q[384]
  PIN i_data_q[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.7850 0.0000 913.8350 0.2200 ;
    END
  END i_data_q[383]
  PIN i_data_q[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.5850 0.0000 913.6350 0.2200 ;
    END
  END i_data_q[382]
  PIN i_data_q[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.3850 0.0000 913.4350 0.2200 ;
    END
  END i_data_q[381]
  PIN i_data_q[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 913.1850 0.0000 913.2350 0.2200 ;
    END
  END i_data_q[380]
  PIN i_data_q[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.7850 0.0000 912.8350 0.2200 ;
    END
  END i_data_q[379]
  PIN i_data_q[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.5850 0.0000 912.6350 0.2200 ;
    END
  END i_data_q[378]
  PIN i_data_q[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.3850 0.0000 912.4350 0.2200 ;
    END
  END i_data_q[377]
  PIN i_data_q[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.1850 0.0000 912.2350 0.2200 ;
    END
  END i_data_q[376]
  PIN i_data_q[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.9850 0.0000 912.0350 0.2200 ;
    END
  END i_data_q[375]
  PIN i_data_q[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.7850 0.0000 911.8350 0.2200 ;
    END
  END i_data_q[374]
  PIN i_data_q[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.5850 0.0000 911.6350 0.2200 ;
    END
  END i_data_q[373]
  PIN i_data_q[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.3850 0.0000 911.4350 0.2200 ;
    END
  END i_data_q[372]
  PIN i_data_q[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 911.1850 0.0000 911.2350 0.2200 ;
    END
  END i_data_q[371]
  PIN i_data_q[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.9850 0.0000 911.0350 0.2200 ;
    END
  END i_data_q[370]
  PIN i_data_q[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.5850 0.0000 910.6350 0.2200 ;
    END
  END i_data_q[369]
  PIN i_data_q[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.3850 0.0000 910.4350 0.2200 ;
    END
  END i_data_q[368]
  PIN i_data_q[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.1850 0.0000 910.2350 0.2200 ;
    END
  END i_data_q[367]
  PIN i_data_q[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.9850 0.0000 910.0350 0.2200 ;
    END
  END i_data_q[366]
  PIN i_data_q[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.7850 0.0000 909.8350 0.2200 ;
    END
  END i_data_q[365]
  PIN i_data_q[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.5850 0.0000 909.6350 0.2200 ;
    END
  END i_data_q[364]
  PIN i_data_q[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.3850 0.0000 909.4350 0.2200 ;
    END
  END i_data_q[363]
  PIN i_data_q[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 909.1850 0.0000 909.2350 0.2200 ;
    END
  END i_data_q[362]
  PIN i_data_q[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.9850 0.0000 909.0350 0.2200 ;
    END
  END i_data_q[361]
  PIN i_data_q[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.7850 0.0000 908.8350 0.2200 ;
    END
  END i_data_q[360]
  PIN i_data_q[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.3850 0.0000 908.4350 0.2200 ;
    END
  END i_data_q[359]
  PIN i_data_q[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.1850 0.0000 908.2350 0.2200 ;
    END
  END i_data_q[358]
  PIN i_data_q[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.9850 0.0000 908.0350 0.2200 ;
    END
  END i_data_q[357]
  PIN i_data_q[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.7850 0.0000 907.8350 0.2200 ;
    END
  END i_data_q[356]
  PIN i_data_q[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.5850 0.0000 907.6350 0.2200 ;
    END
  END i_data_q[355]
  PIN i_data_q[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.3850 0.0000 907.4350 0.2200 ;
    END
  END i_data_q[354]
  PIN i_data_q[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 907.1850 0.0000 907.2350 0.2200 ;
    END
  END i_data_q[353]
  PIN i_data_q[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.9850 0.0000 907.0350 0.2200 ;
    END
  END i_data_q[352]
  PIN i_data_q[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.7850 0.0000 906.8350 0.2200 ;
    END
  END i_data_q[351]
  PIN i_data_q[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.5850 0.0000 906.6350 0.2200 ;
    END
  END i_data_q[350]
  PIN i_data_q[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.1850 0.0000 906.2350 0.2200 ;
    END
  END i_data_q[349]
  PIN i_data_q[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.9850 0.0000 906.0350 0.2200 ;
    END
  END i_data_q[348]
  PIN i_data_q[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.7850 0.0000 905.8350 0.2200 ;
    END
  END i_data_q[347]
  PIN i_data_q[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.5850 0.0000 905.6350 0.2200 ;
    END
  END i_data_q[346]
  PIN i_data_q[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.3850 0.0000 905.4350 0.2200 ;
    END
  END i_data_q[345]
  PIN i_data_q[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 905.1850 0.0000 905.2350 0.2200 ;
    END
  END i_data_q[344]
  PIN i_data_q[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.9850 0.0000 905.0350 0.2200 ;
    END
  END i_data_q[343]
  PIN i_data_q[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.7850 0.0000 904.8350 0.2200 ;
    END
  END i_data_q[342]
  PIN i_data_q[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.5850 0.0000 904.6350 0.2200 ;
    END
  END i_data_q[341]
  PIN i_data_q[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.3850 0.0000 904.4350 0.2200 ;
    END
  END i_data_q[340]
  PIN i_data_q[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.9850 0.0000 904.0350 0.2200 ;
    END
  END i_data_q[339]
  PIN i_data_q[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.7850 0.0000 903.8350 0.2200 ;
    END
  END i_data_q[338]
  PIN i_data_q[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.5850 0.0000 903.6350 0.2200 ;
    END
  END i_data_q[337]
  PIN i_data_q[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.3850 0.0000 903.4350 0.2200 ;
    END
  END i_data_q[336]
  PIN i_data_q[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 903.1850 0.0000 903.2350 0.2200 ;
    END
  END i_data_q[335]
  PIN i_data_q[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.9850 0.0000 903.0350 0.2200 ;
    END
  END i_data_q[334]
  PIN i_data_q[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.7850 0.0000 902.8350 0.2200 ;
    END
  END i_data_q[333]
  PIN i_data_q[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.5850 0.0000 902.6350 0.2200 ;
    END
  END i_data_q[332]
  PIN i_data_q[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.3850 0.0000 902.4350 0.2200 ;
    END
  END i_data_q[331]
  PIN i_data_q[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 902.1850 0.0000 902.2350 0.2200 ;
    END
  END i_data_q[330]
  PIN i_data_q[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 898.1850 0.0000 898.2350 0.2200 ;
    END
  END i_data_q[329]
  PIN i_data_q[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.9850 0.0000 898.0350 0.2200 ;
    END
  END i_data_q[328]
  PIN i_data_q[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.7850 0.0000 897.8350 0.2200 ;
    END
  END i_data_q[327]
  PIN i_data_q[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.5850 0.0000 897.6350 0.2200 ;
    END
  END i_data_q[326]
  PIN i_data_q[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.3850 0.0000 897.4350 0.2200 ;
    END
  END i_data_q[325]
  PIN i_data_q[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 897.1850 0.0000 897.2350 0.2200 ;
    END
  END i_data_q[324]
  PIN i_data_q[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.9850 0.0000 897.0350 0.2200 ;
    END
  END i_data_q[323]
  PIN i_data_q[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.7850 0.0000 896.8350 0.2200 ;
    END
  END i_data_q[322]
  PIN i_data_q[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.5850 0.0000 896.6350 0.2200 ;
    END
  END i_data_q[321]
  PIN i_data_q[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.3850 0.0000 896.4350 0.2200 ;
    END
  END i_data_q[320]
  PIN i_data_q[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.9850 0.0000 896.0350 0.2200 ;
    END
  END i_data_q[319]
  PIN i_data_q[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.7850 0.0000 895.8350 0.2200 ;
    END
  END i_data_q[318]
  PIN i_data_q[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.5850 0.0000 895.6350 0.2200 ;
    END
  END i_data_q[317]
  PIN i_data_q[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.3850 0.0000 895.4350 0.2200 ;
    END
  END i_data_q[316]
  PIN i_data_q[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 895.1850 0.0000 895.2350 0.2200 ;
    END
  END i_data_q[315]
  PIN i_data_q[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.9850 0.0000 895.0350 0.2200 ;
    END
  END i_data_q[314]
  PIN i_data_q[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.7850 0.0000 894.8350 0.2200 ;
    END
  END i_data_q[313]
  PIN i_data_q[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.5850 0.0000 894.6350 0.2200 ;
    END
  END i_data_q[312]
  PIN i_data_q[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.3850 0.0000 894.4350 0.2200 ;
    END
  END i_data_q[311]
  PIN i_data_q[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 894.1850 0.0000 894.2350 0.2200 ;
    END
  END i_data_q[310]
  PIN i_data_q[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.7850 0.0000 893.8350 0.2200 ;
    END
  END i_data_q[309]
  PIN i_data_q[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.5850 0.0000 893.6350 0.2200 ;
    END
  END i_data_q[308]
  PIN i_data_q[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.3850 0.0000 893.4350 0.2200 ;
    END
  END i_data_q[307]
  PIN i_data_q[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.1850 0.0000 893.2350 0.2200 ;
    END
  END i_data_q[306]
  PIN i_data_q[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.9850 0.0000 893.0350 0.2200 ;
    END
  END i_data_q[305]
  PIN i_data_q[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.7850 0.0000 892.8350 0.2200 ;
    END
  END i_data_q[304]
  PIN i_data_q[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.5850 0.0000 892.6350 0.2200 ;
    END
  END i_data_q[303]
  PIN i_data_q[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.3850 0.0000 892.4350 0.2200 ;
    END
  END i_data_q[302]
  PIN i_data_q[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 892.1850 0.0000 892.2350 0.2200 ;
    END
  END i_data_q[301]
  PIN i_data_q[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.9850 0.0000 892.0350 0.2200 ;
    END
  END i_data_q[300]
  PIN i_data_q[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.3850 0.0000 891.4350 0.2200 ;
    END
  END i_data_q[299]
  PIN i_data_q[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.1850 0.0000 891.2350 0.2200 ;
    END
  END i_data_q[298]
  PIN i_data_q[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.9850 0.0000 891.0350 0.2200 ;
    END
  END i_data_q[297]
  PIN i_data_q[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.7850 0.0000 890.8350 0.2200 ;
    END
  END i_data_q[296]
  PIN i_data_q[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.5850 0.0000 890.6350 0.2200 ;
    END
  END i_data_q[295]
  PIN i_data_q[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.3850 0.0000 890.4350 0.2200 ;
    END
  END i_data_q[294]
  PIN i_data_q[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 890.1850 0.0000 890.2350 0.2200 ;
    END
  END i_data_q[293]
  PIN i_data_q[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.9850 0.0000 890.0350 0.2200 ;
    END
  END i_data_q[292]
  PIN i_data_q[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.7850 0.0000 889.8350 0.2200 ;
    END
  END i_data_q[291]
  PIN i_data_q[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.5850 0.0000 889.6350 0.2200 ;
    END
  END i_data_q[290]
  PIN i_data_q[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.1850 0.0000 889.2350 0.2200 ;
    END
  END i_data_q[289]
  PIN i_data_q[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.9850 0.0000 889.0350 0.2200 ;
    END
  END i_data_q[288]
  PIN i_data_q[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.7850 0.0000 888.8350 0.2200 ;
    END
  END i_data_q[287]
  PIN i_data_q[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.5850 0.0000 888.6350 0.2200 ;
    END
  END i_data_q[286]
  PIN i_data_q[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.3850 0.0000 888.4350 0.2200 ;
    END
  END i_data_q[285]
  PIN i_data_q[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 888.1850 0.0000 888.2350 0.2200 ;
    END
  END i_data_q[284]
  PIN i_data_q[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.9850 0.0000 888.0350 0.2200 ;
    END
  END i_data_q[283]
  PIN i_data_q[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.7850 0.0000 887.8350 0.2200 ;
    END
  END i_data_q[282]
  PIN i_data_q[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.5850 0.0000 887.6350 0.2200 ;
    END
  END i_data_q[281]
  PIN i_data_q[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.3850 0.0000 887.4350 0.2200 ;
    END
  END i_data_q[280]
  PIN i_data_q[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.9850 0.0000 887.0350 0.2200 ;
    END
  END i_data_q[279]
  PIN i_data_q[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.7850 0.0000 886.8350 0.2200 ;
    END
  END i_data_q[278]
  PIN i_data_q[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.5850 0.0000 886.6350 0.2200 ;
    END
  END i_data_q[277]
  PIN i_data_q[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.3850 0.0000 886.4350 0.2200 ;
    END
  END i_data_q[276]
  PIN i_data_q[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 886.1850 0.0000 886.2350 0.2200 ;
    END
  END i_data_q[275]
  PIN i_data_q[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.9850 0.0000 886.0350 0.2200 ;
    END
  END i_data_q[274]
  PIN i_data_q[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.7850 0.0000 885.8350 0.2200 ;
    END
  END i_data_q[273]
  PIN i_data_q[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.5850 0.0000 885.6350 0.2200 ;
    END
  END i_data_q[272]
  PIN i_data_q[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.3850 0.0000 885.4350 0.2200 ;
    END
  END i_data_q[271]
  PIN i_data_q[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 885.1850 0.0000 885.2350 0.2200 ;
    END
  END i_data_q[270]
  PIN i_data_q[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.7850 0.0000 884.8350 0.2200 ;
    END
  END i_data_q[269]
  PIN i_data_q[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.5850 0.0000 884.6350 0.2200 ;
    END
  END i_data_q[268]
  PIN i_data_q[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.3850 0.0000 884.4350 0.2200 ;
    END
  END i_data_q[267]
  PIN i_data_q[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.1850 0.0000 884.2350 0.2200 ;
    END
  END i_data_q[266]
  PIN i_data_q[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.9850 0.0000 884.0350 0.2200 ;
    END
  END i_data_q[265]
  PIN i_data_q[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.7850 0.0000 883.8350 0.2200 ;
    END
  END i_data_q[264]
  PIN i_data_q[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.5850 0.0000 883.6350 0.2200 ;
    END
  END i_data_q[263]
  PIN i_data_q[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.3850 0.0000 883.4350 0.2200 ;
    END
  END i_data_q[262]
  PIN i_data_q[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 883.1850 0.0000 883.2350 0.2200 ;
    END
  END i_data_q[261]
  PIN i_data_q[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.9850 0.0000 883.0350 0.2200 ;
    END
  END i_data_q[260]
  PIN i_data_q[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.5850 0.0000 882.6350 0.2200 ;
    END
  END i_data_q[259]
  PIN i_data_q[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.3850 0.0000 882.4350 0.2200 ;
    END
  END i_data_q[258]
  PIN i_data_q[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.1850 0.0000 882.2350 0.2200 ;
    END
  END i_data_q[257]
  PIN i_data_q[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.9850 0.0000 882.0350 0.2200 ;
    END
  END i_data_q[256]
  PIN i_data_q[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.7850 0.0000 881.8350 0.2200 ;
    END
  END i_data_q[255]
  PIN i_data_q[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.5850 0.0000 881.6350 0.2200 ;
    END
  END i_data_q[254]
  PIN i_data_q[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.3850 0.0000 881.4350 0.2200 ;
    END
  END i_data_q[253]
  PIN i_data_q[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 881.1850 0.0000 881.2350 0.2200 ;
    END
  END i_data_q[252]
  PIN i_data_q[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.9850 0.0000 881.0350 0.2200 ;
    END
  END i_data_q[251]
  PIN i_data_q[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.7850 0.0000 880.8350 0.2200 ;
    END
  END i_data_q[250]
  PIN i_data_q[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.3850 0.0000 880.4350 0.2200 ;
    END
  END i_data_q[249]
  PIN i_data_q[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.1850 0.0000 880.2350 0.2200 ;
    END
  END i_data_q[248]
  PIN i_data_q[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.9850 0.0000 880.0350 0.2200 ;
    END
  END i_data_q[247]
  PIN i_data_q[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.7850 0.0000 879.8350 0.2200 ;
    END
  END i_data_q[246]
  PIN i_data_q[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.5850 0.0000 879.6350 0.2200 ;
    END
  END i_data_q[245]
  PIN i_data_q[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.3850 0.0000 879.4350 0.2200 ;
    END
  END i_data_q[244]
  PIN i_data_q[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 879.1850 0.0000 879.2350 0.2200 ;
    END
  END i_data_q[243]
  PIN i_data_q[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.9850 0.0000 879.0350 0.2200 ;
    END
  END i_data_q[242]
  PIN i_data_q[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.7850 0.0000 878.8350 0.2200 ;
    END
  END i_data_q[241]
  PIN i_data_q[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.5850 0.0000 878.6350 0.2200 ;
    END
  END i_data_q[240]
  PIN i_data_q[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.1850 0.0000 878.2350 0.2200 ;
    END
  END i_data_q[239]
  PIN i_data_q[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 877.9850 0.0000 878.0350 0.2200 ;
    END
  END i_data_q[238]
  PIN i_data_q[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 877.7850 0.0000 877.8350 0.2200 ;
    END
  END i_data_q[237]
  PIN i_data_q[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 874.0850 0.0000 874.1350 0.2200 ;
    END
  END i_data_q[236]
  PIN i_data_q[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.8850 0.0000 873.9350 0.2200 ;
    END
  END i_data_q[235]
  PIN i_data_q[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.6850 0.0000 873.7350 0.2200 ;
    END
  END i_data_q[234]
  PIN i_data_q[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.4850 0.0000 873.5350 0.2200 ;
    END
  END i_data_q[233]
  PIN i_data_q[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.2850 0.0000 873.3350 0.2200 ;
    END
  END i_data_q[232]
  PIN i_data_q[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 873.0850 0.0000 873.1350 0.2200 ;
    END
  END i_data_q[231]
  PIN i_data_q[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.8850 0.0000 872.9350 0.2200 ;
    END
  END i_data_q[230]
  PIN i_data_q[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.4850 0.0000 872.5350 0.2200 ;
    END
  END i_data_q[229]
  PIN i_data_q[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.2850 0.0000 872.3350 0.2200 ;
    END
  END i_data_q[228]
  PIN i_data_q[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.0850 0.0000 872.1350 0.2200 ;
    END
  END i_data_q[227]
  PIN i_data_q[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.8850 0.0000 871.9350 0.2200 ;
    END
  END i_data_q[226]
  PIN i_data_q[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.6850 0.0000 871.7350 0.2200 ;
    END
  END i_data_q[225]
  PIN i_data_q[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.4850 0.0000 871.5350 0.2200 ;
    END
  END i_data_q[224]
  PIN i_data_q[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.2850 0.0000 871.3350 0.2200 ;
    END
  END i_data_q[223]
  PIN i_data_q[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 871.0850 0.0000 871.1350 0.2200 ;
    END
  END i_data_q[222]
  PIN i_data_q[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.8850 0.0000 870.9350 0.2200 ;
    END
  END i_data_q[221]
  PIN i_data_q[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.6850 0.0000 870.7350 0.2200 ;
    END
  END i_data_q[220]
  PIN i_data_q[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.2850 0.0000 870.3350 0.2200 ;
    END
  END i_data_q[219]
  PIN i_data_q[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.0850 0.0000 870.1350 0.2200 ;
    END
  END i_data_q[218]
  PIN i_data_q[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.8850 0.0000 869.9350 0.2200 ;
    END
  END i_data_q[217]
  PIN i_data_q[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.6850 0.0000 869.7350 0.2200 ;
    END
  END i_data_q[216]
  PIN i_data_q[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.4850 0.0000 869.5350 0.2200 ;
    END
  END i_data_q[215]
  PIN i_data_q[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.2850 0.0000 869.3350 0.2200 ;
    END
  END i_data_q[214]
  PIN i_data_q[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 869.0850 0.0000 869.1350 0.2200 ;
    END
  END i_data_q[213]
  PIN i_data_q[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.8850 0.0000 868.9350 0.2200 ;
    END
  END i_data_q[212]
  PIN i_data_q[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.6850 0.0000 868.7350 0.2200 ;
    END
  END i_data_q[211]
  PIN i_data_q[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.4850 0.0000 868.5350 0.2200 ;
    END
  END i_data_q[210]
  PIN i_data_q[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.0850 0.0000 868.1350 0.2200 ;
    END
  END i_data_q[209]
  PIN i_data_q[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.8850 0.0000 867.9350 0.2200 ;
    END
  END i_data_q[208]
  PIN i_data_q[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.6850 0.0000 867.7350 0.2200 ;
    END
  END i_data_q[207]
  PIN i_data_q[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.4850 0.0000 867.5350 0.2200 ;
    END
  END i_data_q[206]
  PIN i_data_q[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.2850 0.0000 867.3350 0.2200 ;
    END
  END i_data_q[205]
  PIN i_data_q[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 867.0850 0.0000 867.1350 0.2200 ;
    END
  END i_data_q[204]
  PIN i_data_q[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.8850 0.0000 866.9350 0.2200 ;
    END
  END i_data_q[203]
  PIN i_data_q[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.6850 0.0000 866.7350 0.2200 ;
    END
  END i_data_q[202]
  PIN i_data_q[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.4850 0.0000 866.5350 0.2200 ;
    END
  END i_data_q[201]
  PIN i_data_q[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.2850 0.0000 866.3350 0.2200 ;
    END
  END i_data_q[200]
  PIN i_data_q[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.6850 0.0000 865.7350 0.2200 ;
    END
  END i_data_q[199]
  PIN i_data_q[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.4850 0.0000 865.5350 0.2200 ;
    END
  END i_data_q[198]
  PIN i_data_q[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.2850 0.0000 865.3350 0.2200 ;
    END
  END i_data_q[197]
  PIN i_data_q[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.0850 0.0000 865.1350 0.2200 ;
    END
  END i_data_q[196]
  PIN i_data_q[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.8850 0.0000 864.9350 0.2200 ;
    END
  END i_data_q[195]
  PIN i_data_q[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.6850 0.0000 864.7350 0.2200 ;
    END
  END i_data_q[194]
  PIN i_data_q[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.4850 0.0000 864.5350 0.2200 ;
    END
  END i_data_q[193]
  PIN i_data_q[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.2850 0.0000 864.3350 0.2200 ;
    END
  END i_data_q[192]
  PIN i_data_q[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 864.0850 0.0000 864.1350 0.2200 ;
    END
  END i_data_q[191]
  PIN i_data_q[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.8850 0.0000 863.9350 0.2200 ;
    END
  END i_data_q[190]
  PIN i_data_q[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.4850 0.0000 863.5350 0.2200 ;
    END
  END i_data_q[189]
  PIN i_data_q[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.2850 0.0000 863.3350 0.2200 ;
    END
  END i_data_q[188]
  PIN i_data_q[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.0850 0.0000 863.1350 0.2200 ;
    END
  END i_data_q[187]
  PIN i_data_q[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.8850 0.0000 862.9350 0.2200 ;
    END
  END i_data_q[186]
  PIN i_data_q[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.6850 0.0000 862.7350 0.2200 ;
    END
  END i_data_q[185]
  PIN i_data_q[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.4850 0.0000 862.5350 0.2200 ;
    END
  END i_data_q[184]
  PIN i_data_q[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.2850 0.0000 862.3350 0.2200 ;
    END
  END i_data_q[183]
  PIN i_data_q[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 862.0850 0.0000 862.1350 0.2200 ;
    END
  END i_data_q[182]
  PIN i_data_q[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.8850 0.0000 861.9350 0.2200 ;
    END
  END i_data_q[181]
  PIN i_data_q[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.6850 0.0000 861.7350 0.2200 ;
    END
  END i_data_q[180]
  PIN i_data_q[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.2850 0.0000 861.3350 0.2200 ;
    END
  END i_data_q[179]
  PIN i_data_q[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.0850 0.0000 861.1350 0.2200 ;
    END
  END i_data_q[178]
  PIN i_data_q[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.8850 0.0000 860.9350 0.2200 ;
    END
  END i_data_q[177]
  PIN i_data_q[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.6850 0.0000 860.7350 0.2200 ;
    END
  END i_data_q[176]
  PIN i_data_q[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.4850 0.0000 860.5350 0.2200 ;
    END
  END i_data_q[175]
  PIN i_data_q[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.2850 0.0000 860.3350 0.2200 ;
    END
  END i_data_q[174]
  PIN i_data_q[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 860.0850 0.0000 860.1350 0.2200 ;
    END
  END i_data_q[173]
  PIN i_data_q[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.8850 0.0000 859.9350 0.2200 ;
    END
  END i_data_q[172]
  PIN i_data_q[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.6850 0.0000 859.7350 0.2200 ;
    END
  END i_data_q[171]
  PIN i_data_q[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.4850 0.0000 859.5350 0.2200 ;
    END
  END i_data_q[170]
  PIN i_data_q[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.0850 0.0000 859.1350 0.2200 ;
    END
  END i_data_q[169]
  PIN i_data_q[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.8850 0.0000 858.9350 0.2200 ;
    END
  END i_data_q[168]
  PIN i_data_q[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.6850 0.0000 858.7350 0.2200 ;
    END
  END i_data_q[167]
  PIN i_data_q[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.4850 0.0000 858.5350 0.2200 ;
    END
  END i_data_q[166]
  PIN i_data_q[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.2850 0.0000 858.3350 0.2200 ;
    END
  END i_data_q[165]
  PIN i_data_q[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 858.0850 0.0000 858.1350 0.2200 ;
    END
  END i_data_q[164]
  PIN i_data_q[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.8850 0.0000 857.9350 0.2200 ;
    END
  END i_data_q[163]
  PIN i_data_q[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.6850 0.0000 857.7350 0.2200 ;
    END
  END i_data_q[162]
  PIN i_data_q[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.4850 0.0000 857.5350 0.2200 ;
    END
  END i_data_q[161]
  PIN i_data_q[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.2850 0.0000 857.3350 0.2200 ;
    END
  END i_data_q[160]
  PIN i_data_q[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.8850 0.0000 856.9350 0.2200 ;
    END
  END i_data_q[159]
  PIN i_data_q[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.6850 0.0000 856.7350 0.2200 ;
    END
  END i_data_q[158]
  PIN i_data_q[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.4850 0.0000 856.5350 0.2200 ;
    END
  END i_data_q[157]
  PIN i_data_q[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.2850 0.0000 856.3350 0.2200 ;
    END
  END i_data_q[156]
  PIN i_data_q[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 856.0850 0.0000 856.1350 0.2200 ;
    END
  END i_data_q[155]
  PIN i_data_q[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.8850 0.0000 855.9350 0.2200 ;
    END
  END i_data_q[154]
  PIN i_data_q[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.6850 0.0000 855.7350 0.2200 ;
    END
  END i_data_q[153]
  PIN i_data_q[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.4850 0.0000 855.5350 0.2200 ;
    END
  END i_data_q[152]
  PIN i_data_q[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.2850 0.0000 855.3350 0.2200 ;
    END
  END i_data_q[151]
  PIN i_data_q[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 855.0850 0.0000 855.1350 0.2200 ;
    END
  END i_data_q[150]
  PIN i_data_q[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.6850 0.0000 854.7350 0.2200 ;
    END
  END i_data_q[149]
  PIN i_data_q[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.4850 0.0000 854.5350 0.2200 ;
    END
  END i_data_q[148]
  PIN i_data_q[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.2850 0.0000 854.3350 0.2200 ;
    END
  END i_data_q[147]
  PIN i_data_q[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.0850 0.0000 854.1350 0.2200 ;
    END
  END i_data_q[146]
  PIN i_data_q[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.8850 0.0000 853.9350 0.2200 ;
    END
  END i_data_q[145]
  PIN i_data_q[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.6850 0.0000 853.7350 0.2200 ;
    END
  END i_data_q[144]
  PIN i_data_q[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 853.4850 0.0000 853.5350 0.2200 ;
    END
  END i_data_q[143]
  PIN i_data_q[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.7850 0.0000 849.8350 0.2200 ;
    END
  END i_data_q[142]
  PIN i_data_q[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.5850 0.0000 849.6350 0.2200 ;
    END
  END i_data_q[141]
  PIN i_data_q[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.3850 0.0000 849.4350 0.2200 ;
    END
  END i_data_q[140]
  PIN i_data_q[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.9850 0.0000 849.0350 0.2200 ;
    END
  END i_data_q[139]
  PIN i_data_q[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.7850 0.0000 848.8350 0.2200 ;
    END
  END i_data_q[138]
  PIN i_data_q[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.5850 0.0000 848.6350 0.2200 ;
    END
  END i_data_q[137]
  PIN i_data_q[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.3850 0.0000 848.4350 0.2200 ;
    END
  END i_data_q[136]
  PIN i_data_q[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 848.1850 0.0000 848.2350 0.2200 ;
    END
  END i_data_q[135]
  PIN i_data_q[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.9850 0.0000 848.0350 0.2200 ;
    END
  END i_data_q[134]
  PIN i_data_q[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.7850 0.0000 847.8350 0.2200 ;
    END
  END i_data_q[133]
  PIN i_data_q[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.5850 0.0000 847.6350 0.2200 ;
    END
  END i_data_q[132]
  PIN i_data_q[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.3850 0.0000 847.4350 0.2200 ;
    END
  END i_data_q[131]
  PIN i_data_q[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 847.1850 0.0000 847.2350 0.2200 ;
    END
  END i_data_q[130]
  PIN i_data_q[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.7850 0.0000 846.8350 0.2200 ;
    END
  END i_data_q[129]
  PIN i_data_q[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.5850 0.0000 846.6350 0.2200 ;
    END
  END i_data_q[128]
  PIN i_data_q[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.3850 0.0000 846.4350 0.2200 ;
    END
  END i_data_q[127]
  PIN i_data_q[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.1850 0.0000 846.2350 0.2200 ;
    END
  END i_data_q[126]
  PIN i_data_q[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.9850 0.0000 846.0350 0.2200 ;
    END
  END i_data_q[125]
  PIN i_data_q[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.7850 0.0000 845.8350 0.2200 ;
    END
  END i_data_q[124]
  PIN i_data_q[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.5850 0.0000 845.6350 0.2200 ;
    END
  END i_data_q[123]
  PIN i_data_q[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.3850 0.0000 845.4350 0.2200 ;
    END
  END i_data_q[122]
  PIN i_data_q[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 845.1850 0.0000 845.2350 0.2200 ;
    END
  END i_data_q[121]
  PIN i_data_q[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.9850 0.0000 845.0350 0.2200 ;
    END
  END i_data_q[120]
  PIN i_data_q[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.5850 0.0000 844.6350 0.2200 ;
    END
  END i_data_q[119]
  PIN i_data_q[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.3850 0.0000 844.4350 0.2200 ;
    END
  END i_data_q[118]
  PIN i_data_q[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.1850 0.0000 844.2350 0.2200 ;
    END
  END i_data_q[117]
  PIN i_data_q[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.9850 0.0000 844.0350 0.2200 ;
    END
  END i_data_q[116]
  PIN i_data_q[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.7850 0.0000 843.8350 0.2200 ;
    END
  END i_data_q[115]
  PIN i_data_q[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.5850 0.0000 843.6350 0.2200 ;
    END
  END i_data_q[114]
  PIN i_data_q[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.3850 0.0000 843.4350 0.2200 ;
    END
  END i_data_q[113]
  PIN i_data_q[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 843.1850 0.0000 843.2350 0.2200 ;
    END
  END i_data_q[112]
  PIN i_data_q[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.9850 0.0000 843.0350 0.2200 ;
    END
  END i_data_q[111]
  PIN i_data_q[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.7850 0.0000 842.8350 0.2200 ;
    END
  END i_data_q[110]
  PIN i_data_q[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.3850 0.0000 842.4350 0.2200 ;
    END
  END i_data_q[109]
  PIN i_data_q[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.1850 0.0000 842.2350 0.2200 ;
    END
  END i_data_q[108]
  PIN i_data_q[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.9850 0.0000 842.0350 0.2200 ;
    END
  END i_data_q[107]
  PIN i_data_q[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.7850 0.0000 841.8350 0.2200 ;
    END
  END i_data_q[106]
  PIN i_data_q[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.5850 0.0000 841.6350 0.2200 ;
    END
  END i_data_q[105]
  PIN i_data_q[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.3850 0.0000 841.4350 0.2200 ;
    END
  END i_data_q[104]
  PIN i_data_q[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 841.1850 0.0000 841.2350 0.2200 ;
    END
  END i_data_q[103]
  PIN i_data_q[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.9850 0.0000 841.0350 0.2200 ;
    END
  END i_data_q[102]
  PIN i_data_q[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.7850 0.0000 840.8350 0.2200 ;
    END
  END i_data_q[101]
  PIN i_data_q[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.5850 0.0000 840.6350 0.2200 ;
    END
  END i_data_q[100]
  PIN i_data_q[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.5850 0.0000 976.6350 0.2200 ;
    END
  END i_data_q[99]
  PIN i_data_q[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.3850 0.0000 976.4350 0.2200 ;
    END
  END i_data_q[98]
  PIN i_data_q[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.1850 0.0000 976.2350 0.2200 ;
    END
  END i_data_q[97]
  PIN i_data_q[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.9850 0.0000 976.0350 0.2200 ;
    END
  END i_data_q[96]
  PIN i_data_q[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.7850 0.0000 975.8350 0.2200 ;
    END
  END i_data_q[95]
  PIN i_data_q[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.5850 0.0000 975.6350 0.2200 ;
    END
  END i_data_q[94]
  PIN i_data_q[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.3850 0.0000 975.4350 0.2200 ;
    END
  END i_data_q[93]
  PIN i_data_q[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 975.1850 0.0000 975.2350 0.2200 ;
    END
  END i_data_q[92]
  PIN i_data_q[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.9850 0.0000 975.0350 0.2200 ;
    END
  END i_data_q[91]
  PIN i_data_q[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.7850 0.0000 974.8350 0.2200 ;
    END
  END i_data_q[90]
  PIN i_data_q[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.3850 0.0000 974.4350 0.2200 ;
    END
  END i_data_q[89]
  PIN i_data_q[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.1850 0.0000 974.2350 0.2200 ;
    END
  END i_data_q[88]
  PIN i_data_q[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 970.3850 0.0000 970.4350 0.2200 ;
    END
  END i_data_q[87]
  PIN i_data_q[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 970.1850 0.0000 970.2350 0.2200 ;
    END
  END i_data_q[86]
  PIN i_data_q[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.9850 0.0000 970.0350 0.2200 ;
    END
  END i_data_q[85]
  PIN i_data_q[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.7850 0.0000 969.8350 0.2200 ;
    END
  END i_data_q[84]
  PIN i_data_q[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.5850 0.0000 969.6350 0.2200 ;
    END
  END i_data_q[83]
  PIN i_data_q[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.3850 0.0000 969.4350 0.2200 ;
    END
  END i_data_q[82]
  PIN i_data_q[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 969.1850 0.0000 969.2350 0.2200 ;
    END
  END i_data_q[81]
  PIN i_data_q[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.9850 0.0000 969.0350 0.2200 ;
    END
  END i_data_q[80]
  PIN i_data_q[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.5850 0.0000 968.6350 0.2200 ;
    END
  END i_data_q[79]
  PIN i_data_q[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.3850 0.0000 968.4350 0.2200 ;
    END
  END i_data_q[78]
  PIN i_data_q[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.1850 0.0000 968.2350 0.2200 ;
    END
  END i_data_q[77]
  PIN i_data_q[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.9850 0.0000 968.0350 0.2200 ;
    END
  END i_data_q[76]
  PIN i_data_q[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.7850 0.0000 967.8350 0.2200 ;
    END
  END i_data_q[75]
  PIN i_data_q[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.5850 0.0000 967.6350 0.2200 ;
    END
  END i_data_q[74]
  PIN i_data_q[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.3850 0.0000 967.4350 0.2200 ;
    END
  END i_data_q[73]
  PIN i_data_q[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 967.1850 0.0000 967.2350 0.2200 ;
    END
  END i_data_q[72]
  PIN i_data_q[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.9850 0.0000 967.0350 0.2200 ;
    END
  END i_data_q[71]
  PIN i_data_q[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.7850 0.0000 966.8350 0.2200 ;
    END
  END i_data_q[70]
  PIN i_data_q[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.3850 0.0000 966.4350 0.2200 ;
    END
  END i_data_q[69]
  PIN i_data_q[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.1850 0.0000 966.2350 0.2200 ;
    END
  END i_data_q[68]
  PIN i_data_q[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.9850 0.0000 966.0350 0.2200 ;
    END
  END i_data_q[67]
  PIN i_data_q[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.7850 0.0000 965.8350 0.2200 ;
    END
  END i_data_q[66]
  PIN i_data_q[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.5850 0.0000 965.6350 0.2200 ;
    END
  END i_data_q[65]
  PIN i_data_q[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.3850 0.0000 965.4350 0.2200 ;
    END
  END i_data_q[64]
  PIN i_data_q[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 965.1850 0.0000 965.2350 0.2200 ;
    END
  END i_data_q[63]
  PIN i_data_q[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.9850 0.0000 965.0350 0.2200 ;
    END
  END i_data_q[62]
  PIN i_data_q[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.7850 0.0000 964.8350 0.2200 ;
    END
  END i_data_q[61]
  PIN i_data_q[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.5850 0.0000 964.6350 0.2200 ;
    END
  END i_data_q[60]
  PIN i_data_q[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.1850 0.0000 964.2350 0.2200 ;
    END
  END i_data_q[59]
  PIN i_data_q[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.9850 0.0000 964.0350 0.2200 ;
    END
  END i_data_q[58]
  PIN i_data_q[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 963.7850 0.0000 963.8350 0.2200 ;
    END
  END i_data_q[57]
  PIN i_data_q[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 962.3850 0.0000 962.4350 0.2200 ;
    END
  END i_data_q[56]
  PIN i_data_q[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 960.1850 0.0000 960.2350 0.2200 ;
    END
  END i_data_q[55]
  PIN i_data_q[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 957.9850 0.0000 958.0350 0.2200 ;
    END
  END i_data_q[54]
  PIN i_data_q[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 955.7850 0.0000 955.8350 0.2200 ;
    END
  END i_data_q[53]
  PIN i_data_q[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 953.5850 0.0000 953.6350 0.2200 ;
    END
  END i_data_q[52]
  PIN i_data_q[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 951.3850 0.0000 951.4350 0.2200 ;
    END
  END i_data_q[51]
  PIN i_data_q[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 945.5850 0.0000 945.6350 0.2200 ;
    END
  END i_data_q[50]
  PIN i_data_q[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.1850 0.0000 943.2350 0.2200 ;
    END
  END i_data_q[49]
  PIN i_data_q[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 940.9850 0.0000 941.0350 0.2200 ;
    END
  END i_data_q[48]
  PIN i_data_q[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 938.7850 0.0000 938.8350 0.2200 ;
    END
  END i_data_q[47]
  PIN i_data_q[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 936.5850 0.0000 936.6350 0.2200 ;
    END
  END i_data_q[46]
  PIN i_data_q[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 934.3850 0.0000 934.4350 0.2200 ;
    END
  END i_data_q[45]
  PIN i_data_q[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 932.1850 0.0000 932.2350 0.2200 ;
    END
  END i_data_q[44]
  PIN i_data_q[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 929.9850 0.0000 930.0350 0.2200 ;
    END
  END i_data_q[43]
  PIN i_data_q[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 927.7850 0.0000 927.8350 0.2200 ;
    END
  END i_data_q[42]
  PIN i_data_q[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 921.9850 0.0000 922.0350 0.2200 ;
    END
  END i_data_q[41]
  PIN i_data_q[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 919.7850 0.0000 919.8350 0.2200 ;
    END
  END i_data_q[40]
  PIN i_data_q[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.3850 0.0000 917.4350 0.2200 ;
    END
  END i_data_q[39]
  PIN i_data_q[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 915.1850 0.0000 915.2350 0.2200 ;
    END
  END i_data_q[38]
  PIN i_data_q[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 912.9850 0.0000 913.0350 0.2200 ;
    END
  END i_data_q[37]
  PIN i_data_q[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 910.7850 0.0000 910.8350 0.2200 ;
    END
  END i_data_q[36]
  PIN i_data_q[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 908.5850 0.0000 908.6350 0.2200 ;
    END
  END i_data_q[35]
  PIN i_data_q[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 906.3850 0.0000 906.4350 0.2200 ;
    END
  END i_data_q[34]
  PIN i_data_q[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 904.1850 0.0000 904.2350 0.2200 ;
    END
  END i_data_q[33]
  PIN i_data_q[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 898.3850 0.0000 898.4350 0.2200 ;
    END
  END i_data_q[32]
  PIN i_data_q[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 896.1850 0.0000 896.2350 0.2200 ;
    END
  END i_data_q[31]
  PIN i_data_q[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 893.9850 0.0000 894.0350 0.2200 ;
    END
  END i_data_q[30]
  PIN i_data_q[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.5850 0.0000 891.6350 0.2200 ;
    END
  END i_data_q[29]
  PIN i_data_q[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 889.3850 0.0000 889.4350 0.2200 ;
    END
  END i_data_q[28]
  PIN i_data_q[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 887.1850 0.0000 887.2350 0.2200 ;
    END
  END i_data_q[27]
  PIN i_data_q[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 884.9850 0.0000 885.0350 0.2200 ;
    END
  END i_data_q[26]
  PIN i_data_q[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 882.7850 0.0000 882.8350 0.2200 ;
    END
  END i_data_q[25]
  PIN i_data_q[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 880.5850 0.0000 880.6350 0.2200 ;
    END
  END i_data_q[24]
  PIN i_data_q[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 878.3850 0.0000 878.4350 0.2200 ;
    END
  END i_data_q[23]
  PIN i_data_q[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 872.6850 0.0000 872.7350 0.2200 ;
    END
  END i_data_q[22]
  PIN i_data_q[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 870.4850 0.0000 870.5350 0.2200 ;
    END
  END i_data_q[21]
  PIN i_data_q[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 868.2850 0.0000 868.3350 0.2200 ;
    END
  END i_data_q[20]
  PIN i_data_q[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 865.8850 0.0000 865.9350 0.2200 ;
    END
  END i_data_q[19]
  PIN i_data_q[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 863.6850 0.0000 863.7350 0.2200 ;
    END
  END i_data_q[18]
  PIN i_data_q[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 861.4850 0.0000 861.5350 0.2200 ;
    END
  END i_data_q[17]
  PIN i_data_q[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 859.2850 0.0000 859.3350 0.2200 ;
    END
  END i_data_q[16]
  PIN i_data_q[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 857.0850 0.0000 857.1350 0.2200 ;
    END
  END i_data_q[15]
  PIN i_data_q[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 854.8850 0.0000 854.9350 0.2200 ;
    END
  END i_data_q[14]
  PIN i_data_q[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 849.1850 0.0000 849.2350 0.2200 ;
    END
  END i_data_q[13]
  PIN i_data_q[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 846.9850 0.0000 847.0350 0.2200 ;
    END
  END i_data_q[12]
  PIN i_data_q[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 844.7850 0.0000 844.8350 0.2200 ;
    END
  END i_data_q[11]
  PIN i_data_q[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 842.5850 0.0000 842.6350 0.2200 ;
    END
  END i_data_q[10]
  PIN i_data_q[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 976.7850 0.0000 976.8350 0.2200 ;
    END
  END i_data_q[9]
  PIN i_data_q[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 974.5850 0.0000 974.6350 0.2200 ;
    END
  END i_data_q[8]
  PIN i_data_q[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 968.7850 0.0000 968.8350 0.2200 ;
    END
  END i_data_q[7]
  PIN i_data_q[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 966.5850 0.0000 966.6350 0.2200 ;
    END
  END i_data_q[6]
  PIN i_data_q[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 964.3850 0.0000 964.4350 0.2200 ;
    END
  END i_data_q[5]
  PIN i_data_q[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 943.3850 0.0000 943.4350 0.2200 ;
    END
  END i_data_q[4]
  PIN i_data_q[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 917.5850 0.0000 917.6350 0.2200 ;
    END
  END i_data_q[3]
  PIN i_data_q[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 891.7850 0.0000 891.8350 0.2200 ;
    END
  END i_data_q[2]
  PIN i_data_q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 866.0850 0.0000 866.1350 0.2200 ;
    END
  END i_data_q[1]
  PIN i_data_q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 840.3850 0.0000 840.4350 0.2200 ;
    END
  END i_data_q[0]
  PIN i_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1555.8100 0.0000 1555.9100 0.4000 ;
    END
  END i_valid
  PIN o_fo_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.2850 640.5800 1701.3350 640.8000 ;
    END
  END o_fo_valid
  PIN o_fo_value[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.6850 640.5800 1703.7350 640.8000 ;
    END
  END o_fo_value[14]
  PIN o_fo_value[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 159.8250 1704.3000 159.8750 ;
    END
  END o_fo_value[13]
  PIN o_fo_value[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 191.0250 1704.3000 191.0750 ;
    END
  END o_fo_value[12]
  PIN o_fo_value[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 207.8250 1704.3000 207.8750 ;
    END
  END o_fo_value[11]
  PIN o_fo_value[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 160.5250 1704.3000 160.5750 ;
    END
  END o_fo_value[10]
  PIN o_fo_value[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 163.4250 1704.3000 163.4750 ;
    END
  END o_fo_value[9]
  PIN o_fo_value[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.6850 640.5800 1703.7350 640.8000 ;
    END
  END o_fo_value[8]
  PIN o_fo_value[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.4850 640.5800 1703.5350 640.8000 ;
    END
  END o_fo_value[7]
  PIN o_fo_value[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.4850 640.5800 1703.5350 640.8000 ;
    END
  END o_fo_value[6]
  PIN o_fo_value[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.2850 640.5800 1703.3350 640.8000 ;
    END
  END o_fo_value[5]
  PIN o_fo_value[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.2850 640.5800 1703.3350 640.8000 ;
    END
  END o_fo_value[4]
  PIN o_fo_value[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1703.2100 640.4000 1703.3100 640.8000 ;
    END
  END o_fo_value[3]
  PIN o_fo_value[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.0850 640.5800 1703.1350 640.8000 ;
    END
  END o_fo_value[2]
  PIN o_fo_value[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.0850 640.5800 1703.1350 640.8000 ;
    END
  END o_fo_value[1]
  PIN o_fo_value[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.8850 640.5800 1702.9350 640.8000 ;
    END
  END o_fo_value[0]
  PIN i_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 637.8250 1704.3000 637.8750 ;
    END
  END i_enable
  PIN i_subsampling
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.2850 640.5800 1701.3350 640.8000 ;
    END
  END i_subsampling
  PIN i_static_coef[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 640.2250 1704.3000 640.2750 ;
    END
  END i_static_coef[44]
  PIN i_static_coef[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 640.2250 1704.3000 640.2750 ;
    END
  END i_static_coef[43]
  PIN i_static_coef[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 640.0250 1704.3000 640.0750 ;
    END
  END i_static_coef[42]
  PIN i_static_coef[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 640.0250 1704.3000 640.0750 ;
    END
  END i_static_coef[41]
  PIN i_static_coef[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.8250 1704.3000 639.8750 ;
    END
  END i_static_coef[40]
  PIN i_static_coef[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.8250 1704.3000 639.8750 ;
    END
  END i_static_coef[39]
  PIN i_static_coef[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.6250 1704.3000 639.6750 ;
    END
  END i_static_coef[38]
  PIN i_static_coef[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.6250 1704.3000 639.6750 ;
    END
  END i_static_coef[37]
  PIN i_static_coef[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.4250 1704.3000 639.4750 ;
    END
  END i_static_coef[36]
  PIN i_static_coef[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.4250 1704.3000 639.4750 ;
    END
  END i_static_coef[35]
  PIN i_static_coef[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.8850 640.5800 1702.9350 640.8000 ;
    END
  END i_static_coef[34]
  PIN i_static_coef[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.8100 640.4000 1702.9100 640.8000 ;
    END
  END i_static_coef[33]
  PIN i_static_coef[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.2250 1704.3000 639.2750 ;
    END
  END i_static_coef[32]
  PIN i_static_coef[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.2250 1704.3000 639.2750 ;
    END
  END i_static_coef[31]
  PIN i_static_coef[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.6850 640.5800 1702.7350 640.8000 ;
    END
  END i_static_coef[30]
  PIN i_static_coef[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.6850 640.5800 1702.7350 640.8000 ;
    END
  END i_static_coef[29]
  PIN i_static_coef[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 639.0250 1704.3000 639.0750 ;
    END
  END i_static_coef[28]
  PIN i_static_coef[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 639.0250 1704.3000 639.0750 ;
    END
  END i_static_coef[27]
  PIN i_static_coef[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.4850 640.5800 1702.5350 640.8000 ;
    END
  END i_static_coef[26]
  PIN i_static_coef[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.4850 640.5800 1702.5350 640.8000 ;
    END
  END i_static_coef[25]
  PIN i_static_coef[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.4100 640.4000 1702.5100 640.8000 ;
    END
  END i_static_coef[24]
  PIN i_static_coef[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.8250 1704.3000 638.8750 ;
    END
  END i_static_coef[23]
  PIN i_static_coef[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.5250 1704.3000 0.5750 ;
    END
  END i_static_coef[22]
  PIN i_static_coef[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.8250 1704.3000 638.8750 ;
    END
  END i_static_coef[21]
  PIN i_static_coef[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.2850 640.5800 1702.3350 640.8000 ;
    END
  END i_static_coef[20]
  PIN i_static_coef[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.5250 1704.3000 0.5750 ;
    END
  END i_static_coef[19]
  PIN i_static_coef[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.6850 0.0000 1703.7350 0.2200 ;
    END
  END i_static_coef[18]
  PIN i_static_coef[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.2850 640.5800 1702.3350 640.8000 ;
    END
  END i_static_coef[17]
  PIN i_static_coef[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.6250 1704.3000 638.6750 ;
    END
  END i_static_coef[16]
  PIN i_static_coef[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.6850 0.0000 1703.7350 0.2200 ;
    END
  END i_static_coef[15]
  PIN i_static_coef[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.6250 1704.3000 638.6750 ;
    END
  END i_static_coef[14]
  PIN i_static_coef[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.7250 1704.3000 0.7750 ;
    END
  END i_static_coef[13]
  PIN i_static_coef[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.7250 1704.3000 0.7750 ;
    END
  END i_static_coef[12]
  PIN i_static_coef[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.4850 0.0000 1703.5350 0.2200 ;
    END
  END i_static_coef[11]
  PIN i_static_coef[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1703.4850 0.0000 1703.5350 0.2200 ;
    END
  END i_static_coef[10]
  PIN i_static_coef[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1702.0850 640.5800 1702.1350 640.8000 ;
    END
  END i_static_coef[9]
  PIN i_static_coef[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 0.9250 1704.3000 0.9750 ;
    END
  END i_static_coef[8]
  PIN i_static_coef[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 0.9250 1704.3000 0.9750 ;
    END
  END i_static_coef[7]
  PIN i_static_coef[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1702.0850 640.5800 1702.1350 640.8000 ;
    END
  END i_static_coef[6]
  PIN i_static_coef[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1702.0100 640.4000 1702.1100 640.8000 ;
    END
  END i_static_coef[5]
  PIN i_static_coef[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.4250 1704.3000 638.4750 ;
    END
  END i_static_coef[4]
  PIN i_static_coef[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.4250 1704.3000 638.4750 ;
    END
  END i_static_coef[3]
  PIN i_static_coef[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.8850 640.5800 1701.9350 640.8000 ;
    END
  END i_static_coef[2]
  PIN i_static_coef[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.8850 640.5800 1701.9350 640.8000 ;
    END
  END i_static_coef[1]
  PIN i_static_coef[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1703.2850 0.0000 1703.3350 0.2200 ;
    END
  END i_static_coef[0]
  PIN i_static_pipe_lat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.2250 1704.3000 638.2750 ;
    END
  END i_static_pipe_lat[9]
  PIN i_static_pipe_lat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.2250 1704.3000 638.2750 ;
    END
  END i_static_pipe_lat[8]
  PIN i_static_pipe_lat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.6850 640.5800 1701.7350 640.8000 ;
    END
  END i_static_pipe_lat[7]
  PIN i_static_pipe_lat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.6850 640.5800 1701.7350 640.8000 ;
    END
  END i_static_pipe_lat[6]
  PIN i_static_pipe_lat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1701.6100 640.4000 1701.7100 640.8000 ;
    END
  END i_static_pipe_lat[5]
  PIN i_static_pipe_lat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 638.0250 1704.3000 638.0750 ;
    END
  END i_static_pipe_lat[4]
  PIN i_static_pipe_lat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 1704.0800 638.0250 1704.3000 638.0750 ;
    END
  END i_static_pipe_lat[3]
  PIN i_static_pipe_lat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1701.4850 640.5800 1701.5350 640.8000 ;
    END
  END i_static_pipe_lat[2]
  PIN i_static_pipe_lat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 1701.4850 640.5800 1701.5350 640.8000 ;
    END
  END i_static_pipe_lat[1]
  PIN i_static_pipe_lat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 637.8250 1704.3000 637.8750 ;
    END
  END i_static_pipe_lat[0]
  PIN sc_di0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 51.6850 0.0000 51.7350 0.2200 ;
    END
  END sc_di0
  PIN sc_di1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 51.6850 0.0000 51.7350 0.2200 ;
    END
  END sc_di1
  PIN sc_di2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 115.1250 0.2200 115.1750 ;
    END
  END sc_di2
  PIN sc_di3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 272.6250 0.2200 272.6750 ;
    END
  END sc_di3
  PIN sc_di4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 430.1250 0.2200 430.1750 ;
    END
  END sc_di4
  PIN sc_cpren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 3.3250 0.2200 3.3750 ;
    END
  END sc_cpren
  PIN sc_sen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.4850 0.0000 0.5350 0.2200 ;
    END
  END sc_sen
  PIN sc_spren
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 0.0000 1.4250 0.2200 1.4750 ;
    END
  END sc_spren
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER B1 ;
        RECT 1701.2100 640.4000 1701.3100 640.8000 ;
    END
  END clk
  PIN rst_async_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 1704.0800 637.6250 1704.3000 637.6750 ;
    END
  END rst_async_n
  PIN sc_do0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 1.3850 0.0000 1.4350 0.2200 ;
    END
  END sc_do0
  PIN sc_do1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.2850 0.0000 2.3350 0.2200 ;
    END
  END sc_do1
  PIN sc_do2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.7850 0.0000 0.8350 0.2200 ;
    END
  END sc_do2
  PIN sc_do3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 2.6850 0.0000 2.7350 0.2200 ;
    END
  END sc_do3
  PIN sc_do4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 8.4850 0.0000 8.5350 0.2200 ;
    END
  END sc_do4
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER LB ;
        RECT 1696.8600 191.2960 1704.3000 221.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 546.8400 1704.3000 576.8400 ;
    END
    PORT
      LAYER IA ;
        RECT 1439.9020 640.4000 1446.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1415.9020 640.4000 1422.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1319.9020 640.4000 1326.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1343.9020 640.4000 1350.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1367.9020 640.4000 1374.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1391.9020 640.4000 1398.9020 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 546.8400 1726.8600 621.2200 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 553.1330 1704.3000 553.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 550.7330 1704.3000 550.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 548.3330 1704.3000 548.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 545.9330 1704.3000 546.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 543.5330 1704.3000 543.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 541.1330 1704.3000 541.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 538.7330 1704.3000 538.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 536.3330 1704.3000 536.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 533.9330 1704.3000 534.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 531.5330 1704.3000 531.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 529.1330 1704.3000 529.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 526.7330 1704.3000 526.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 1463.9020 534.8400 1704.3000 541.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 524.3330 1704.3000 524.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 521.9330 1704.3000 522.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 519.5330 1704.3000 519.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 517.1330 1704.3000 517.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 514.7330 1704.3000 514.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 512.3330 1704.3000 512.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 509.9330 1704.3000 510.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 507.5330 1704.3000 507.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 1463.9020 510.8400 1704.3000 517.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1443.0160 606.2200 1506.3080 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 191.2960 1726.8600 265.6760 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 197.9330 1704.3000 198.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 195.5330 1704.3000 195.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 193.1330 1704.3000 193.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 190.7330 1704.3000 190.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 188.3330 1704.3000 188.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 185.9330 1704.3000 186.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 183.5330 1704.3000 183.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 1463.9020 179.2960 1704.3000 186.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 181.1330 1704.3000 181.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 178.7330 1704.3000 178.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 176.3330 1704.3000 176.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 173.9330 1704.3000 174.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 171.5330 1704.3000 171.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 169.1330 1704.3000 169.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 166.7330 1704.3000 166.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 164.3330 1704.3000 164.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 161.9330 1704.3000 162.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 159.5330 1704.3000 159.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 157.1330 1704.3000 157.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 154.7330 1704.3000 154.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 152.3330 1704.3000 152.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 1463.9020 155.2960 1704.3000 162.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1443.0160 250.6760 1506.3080 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 1417.4020 531.8400 1447.4020 610.6060 ;
    END
    PORT
      LAYER LB ;
        RECT 1417.4020 176.2960 1447.4020 255.0620 ;
    END
    PORT
      LAYER LB ;
        RECT 1331.9020 531.8400 1361.9020 576.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 546.8400 1361.9020 576.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 546.8400 1315.7560 621.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 191.2960 1315.7560 265.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 1331.9020 176.2960 1361.9020 221.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 191.2960 1361.9020 221.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1052.7980 534.8400 1310.9020 541.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1052.7980 510.8400 1310.9020 517.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1052.7980 179.2960 1310.9020 186.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1052.7980 155.2960 1310.9020 162.2960 ;
    END
    PORT
      LAYER IA ;
        RECT 956.7980 640.4000 963.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 980.7980 640.4000 987.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1004.7980 640.4000 1011.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1028.7980 640.4000 1035.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 932.7980 640.4000 939.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 908.7980 640.4000 915.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 617.6940 640.4000 624.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 497.6940 640.4000 504.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 521.6940 640.4000 528.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 545.6940 640.4000 552.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 569.6940 640.4000 576.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 593.6940 640.4000 600.6940 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1031.9120 606.2200 1095.2040 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 1006.2980 531.8400 1036.2980 610.6060 ;
    END
    PORT
      LAYER LB ;
        RECT 920.7980 531.8400 950.7980 576.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 546.8400 950.7980 576.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 546.8400 904.6520 621.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 1031.9120 250.6760 1095.2040 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 1006.2980 176.2960 1036.2980 255.0620 ;
    END
    PORT
      LAYER LB ;
        RECT 920.7980 176.2960 950.7980 221.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 191.2960 950.7980 221.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 191.2960 904.6520 265.6760 ;
    END
    PORT
      LAYER IB ;
        RECT 641.6940 534.8400 899.7980 541.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 641.6940 510.8400 899.7980 517.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 641.6940 179.2960 899.7980 186.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 641.6940 155.2960 899.7980 162.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 531.8400 625.1940 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 606.2200 670.1000 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 464.5470 606.2200 539.6940 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 509.6940 531.8400 539.6940 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 176.2960 625.1940 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 250.6760 670.1000 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 464.5470 250.6760 539.6940 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 509.6940 176.2960 539.6940 280.6760 ;
    END
    PORT
      LAYER IB ;
        RECT 230.5900 534.8400 488.6940 541.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 230.5900 510.8400 488.6940 517.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 230.5900 179.2960 488.6940 186.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 230.5900 155.2960 488.6940 162.2960 ;
    END
    PORT
      LAYER IA ;
        RECT 134.5900 640.4000 141.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 158.5900 640.4000 165.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 182.5900 640.4000 189.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 206.5900 640.4000 213.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 86.5900 640.4000 93.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 110.5900 640.4000 117.5900 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 606.2200 258.9960 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 531.8400 214.0900 636.2200 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 250.6760 258.9960 280.6760 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 176.2960 214.0900 280.6760 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 553.1330 0.0500 553.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 550.7330 0.0500 550.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 548.3330 0.0500 548.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 545.9330 0.0500 546.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 543.5330 0.0500 543.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 541.1330 0.0500 541.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 538.7330 0.0500 538.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 536.3330 0.0500 536.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 533.9330 0.0500 534.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 531.5330 0.0500 531.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 529.1330 0.0500 529.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 526.7330 0.0500 526.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 524.3330 0.0500 524.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 521.9330 0.0500 522.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 519.5330 0.0500 519.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 517.1330 0.0500 517.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 514.7330 0.0500 514.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 512.3330 0.0500 512.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 509.9330 0.0500 510.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 507.5330 0.0500 507.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 510.8400 77.5900 517.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 534.8400 77.5900 541.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 197.9330 0.0500 198.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 195.5330 0.0500 195.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 193.1330 0.0500 193.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 190.7330 0.0500 190.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 188.3330 0.0500 188.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 185.9330 0.0500 186.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 183.5330 0.0500 183.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 181.1330 0.0500 181.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 178.7330 0.0500 178.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 176.3330 0.0500 176.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 173.9330 0.0500 174.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 171.5330 0.0500 171.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 169.1330 0.0500 169.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 166.7330 0.0500 166.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 164.3330 0.0500 164.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 161.9330 0.0500 162.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 159.5330 0.0500 159.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 157.1330 0.0500 157.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 154.7330 0.0500 154.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 152.3330 0.0500 152.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 155.2960 77.5900 162.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 179.2960 77.5900 186.2960 ;
    END
    PORT
      LAYER IA ;
        RECT 1682.5370 0.0000 1689.5370 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1682.5370 640.4000 1689.5370 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1658.2270 0.0000 1665.2270 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1658.2270 640.4000 1665.2270 640.8000 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 1.1330 1704.3000 1.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 1.1330 0.0500 1.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 3.5330 1704.3000 3.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 3.5330 0.0500 3.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 5.9330 1704.3000 6.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 5.9330 0.0500 6.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 8.3330 1704.3000 8.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 8.3330 0.0500 8.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 10.7330 1704.3000 10.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 10.7330 0.0500 10.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 13.1330 1704.3000 13.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 13.1330 0.0500 13.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 15.5330 1704.3000 15.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 15.5330 0.0500 15.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 13.3340 1704.3000 20.3340 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 17.9330 1704.3000 18.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 17.9330 0.0500 18.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 20.3330 1704.3000 20.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 20.3330 0.0500 20.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 22.7330 1704.3000 22.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 22.7330 0.0500 22.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 25.1330 1704.3000 25.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 25.1330 0.0500 25.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 27.5330 1704.3000 27.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 27.5330 0.0500 27.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 29.9330 1704.3000 30.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 29.9330 0.0500 30.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 32.3330 1704.3000 32.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 32.3330 0.0500 32.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 34.7330 1704.3000 34.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 34.7330 0.0500 34.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 37.1330 1704.3000 37.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 37.1330 0.0500 37.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 39.5330 1704.3000 39.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 39.5330 0.0500 39.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 41.9330 1704.3000 42.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 41.9330 0.0500 42.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 36.9620 1704.3000 43.9620 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 44.3330 1704.3000 44.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 44.3330 0.0500 44.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 46.7330 1704.3000 46.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 46.7330 0.0500 46.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 49.1330 1704.3000 49.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 49.1330 0.0500 49.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 51.5330 1704.3000 51.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 51.5330 0.0500 51.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 53.9330 1704.3000 54.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 53.9330 0.0500 54.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 56.3330 1704.3000 56.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 56.3330 0.0500 56.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 58.7330 1704.3000 58.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 58.7330 0.0500 58.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 61.1330 1704.3000 61.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 61.1330 0.0500 61.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 60.5900 1704.3000 67.5900 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 63.5330 1704.3000 63.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 63.5330 0.0500 63.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 65.9330 1704.3000 66.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 65.9330 0.0500 66.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 68.3330 1704.3000 68.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 68.3330 0.0500 68.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 70.7330 1704.3000 70.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 70.7330 0.0500 70.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 73.1330 1704.3000 73.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 73.1330 0.0500 73.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 75.5330 1704.3000 75.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 75.5330 0.0500 75.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 77.9330 1704.3000 78.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 77.9330 0.0500 78.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 80.3330 1704.3000 80.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 80.3330 0.0500 80.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 82.7330 1704.3000 82.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 82.7330 0.0500 82.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 85.1330 1704.3000 85.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 85.1330 0.0500 85.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 87.5330 1704.3000 87.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 87.5330 0.0500 87.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 84.2180 1704.3000 91.2180 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 89.9330 1704.3000 90.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 89.9330 0.0500 90.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 92.3330 1704.3000 92.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 92.3330 0.0500 92.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 94.7330 1704.3000 94.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 94.7330 0.0500 94.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 97.1330 1704.3000 97.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 97.1330 0.0500 97.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 99.5330 1704.3000 99.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 99.5330 0.0500 99.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 101.9330 1704.3000 102.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 101.9330 0.0500 102.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 104.3330 1704.3000 104.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 104.3330 0.0500 104.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 106.7330 1704.3000 106.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 106.7330 0.0500 106.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 109.1330 1704.3000 109.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 109.1330 0.0500 109.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 111.5330 1704.3000 111.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 111.5330 0.0500 111.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 107.8460 1704.3000 114.8460 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 113.9330 1704.3000 114.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 113.9330 0.0500 114.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 116.3330 1704.3000 116.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 116.3330 0.0500 116.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 118.7330 1704.3000 118.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 118.7330 0.0500 118.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 121.1330 1704.3000 121.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 121.1330 0.0500 121.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 123.5330 1704.3000 123.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 123.5330 0.0500 123.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 125.9330 1704.3000 126.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 125.9330 0.0500 126.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 128.3330 1704.3000 128.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 128.3330 0.0500 128.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 130.7330 1704.3000 130.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 130.7330 0.0500 130.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 133.1330 1704.3000 133.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 133.1330 0.0500 133.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 131.4740 1704.3000 138.4740 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 135.5330 1704.3000 135.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 135.5330 0.0500 135.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 137.9330 1704.3000 138.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 137.9330 0.0500 138.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 142.7330 1704.3000 142.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 142.7330 0.0500 142.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 140.3330 1704.3000 140.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 140.3330 0.0500 140.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 147.5330 1704.3000 147.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 147.5330 0.0500 147.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 145.1330 1704.3000 145.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 145.1330 0.0500 145.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 149.9330 1704.3000 150.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 149.9330 0.0500 150.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 200.3330 1704.3000 200.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 200.3330 0.0500 200.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 202.7330 1704.3000 202.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 202.7330 0.0500 202.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 203.2960 1704.3000 210.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 205.1330 1704.3000 205.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 205.1330 0.0500 205.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 207.5330 1704.3000 207.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 207.5330 0.0500 207.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 212.3330 1704.3000 212.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 212.3330 0.0500 212.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 209.9330 1704.3000 210.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 209.9330 0.0500 210.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 217.1330 1704.3000 217.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 217.1330 0.0500 217.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 214.7330 1704.3000 214.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 214.7330 0.0500 214.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 221.9330 1704.3000 222.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 221.9330 0.0500 222.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 219.5330 1704.3000 219.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 219.5330 0.0500 219.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 226.7330 1704.3000 226.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 226.7330 0.0500 226.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 224.3330 1704.3000 224.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 224.3330 0.0500 224.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 231.5330 1704.3000 231.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 231.5330 0.0500 231.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 229.1330 1704.3000 229.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 229.1330 0.0500 229.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 227.1100 1704.3000 234.1100 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 233.9330 1704.3000 234.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 233.9330 0.0500 234.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 238.7330 1704.3000 238.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 238.7330 0.0500 238.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 236.3330 1704.3000 236.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 236.3330 0.0500 236.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 243.5330 1704.3000 243.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 243.5330 0.0500 243.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 241.1330 1704.3000 241.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 241.1330 0.0500 241.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 248.3330 1704.3000 248.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 248.3330 0.0500 248.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 245.9330 1704.3000 246.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 245.9330 0.0500 246.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 253.1330 1704.3000 253.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 253.1330 0.0500 253.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 250.7330 1704.3000 250.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 250.7330 0.0500 250.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 250.7380 1704.3000 257.7380 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 257.9330 1704.3000 258.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 257.9330 0.0500 258.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 255.5330 1704.3000 255.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 255.5330 0.0500 255.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 260.3330 1704.3000 260.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 260.3330 0.0500 260.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 262.7330 1704.3000 262.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 262.7330 0.0500 262.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 267.5330 1704.3000 267.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 267.5330 0.0500 267.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 265.1330 1704.3000 265.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 265.1330 0.0500 265.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 272.3330 1704.3000 272.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 272.3330 0.0500 272.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 269.9330 1704.3000 270.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 269.9330 0.0500 270.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 277.1330 1704.3000 277.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 277.1330 0.0500 277.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 274.7330 1704.3000 274.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 274.7330 0.0500 274.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 274.3660 1704.3000 281.3660 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 281.9330 1704.3000 282.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 281.9330 0.0500 282.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 279.5330 1704.3000 279.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 279.5330 0.0500 279.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 289.1330 1704.3000 289.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 289.1330 0.0500 289.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 286.7330 1704.3000 286.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 286.7330 0.0500 286.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 284.3330 1704.3000 284.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 284.3330 0.0500 284.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 293.9330 1704.3000 294.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 293.9330 0.0500 294.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 291.5330 1704.3000 291.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 291.5330 0.0500 291.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 298.7330 1704.3000 298.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 298.7330 0.0500 298.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 296.3330 1704.3000 296.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 296.3330 0.0500 296.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 303.5330 1704.3000 303.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 303.5330 0.0500 303.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 301.1330 1704.3000 301.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 301.1330 0.0500 301.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 297.9940 1704.3000 304.9940 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 308.3330 1704.3000 308.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 308.3330 0.0500 308.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 305.9330 1704.3000 306.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 305.9330 0.0500 306.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 313.1330 1704.3000 313.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 313.1330 0.0500 313.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 310.7330 1704.3000 310.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 310.7330 0.0500 310.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 317.9330 1704.3000 318.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 317.9330 0.0500 318.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 315.5330 1704.3000 315.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 315.5330 0.0500 315.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 322.7330 1704.3000 322.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 322.7330 0.0500 322.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 320.3330 1704.3000 320.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 320.3330 0.0500 320.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 321.6220 1704.3000 328.6220 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 327.5330 1704.3000 327.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 327.5330 0.0500 327.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 325.1330 1704.3000 325.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 325.1330 0.0500 325.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 332.3330 1704.3000 332.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 332.3330 0.0500 332.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 329.9330 1704.3000 330.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 329.9330 0.0500 330.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 337.1330 1704.3000 337.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 337.1330 0.0500 337.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 334.7330 1704.3000 334.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 334.7330 0.0500 334.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 339.5330 1704.3000 339.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 339.5330 0.0500 339.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 344.3330 1704.3000 344.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 344.3330 0.0500 344.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 341.9330 1704.3000 342.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 341.9330 0.0500 342.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 349.1330 1704.3000 349.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 349.1330 0.0500 349.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 346.7330 1704.3000 346.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 346.7330 0.0500 346.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 345.2500 1704.3000 352.2500 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 353.9330 1704.3000 354.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 353.9330 0.0500 354.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 351.5330 1704.3000 351.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 351.5330 0.0500 351.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 356.3330 1704.3000 356.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 356.3330 0.0500 356.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 358.7330 1704.3000 358.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 358.7330 0.0500 358.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 363.5330 1704.3000 363.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 363.5330 0.0500 363.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 361.1330 1704.3000 361.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 361.1330 0.0500 361.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 368.3330 1704.3000 368.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 368.3330 0.0500 368.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 365.9330 1704.3000 366.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 365.9330 0.0500 366.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 373.1330 1704.3000 373.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 373.1330 0.0500 373.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 370.7330 1704.3000 370.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 370.7330 0.0500 370.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 368.8780 1704.3000 375.8780 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 375.5330 1704.3000 375.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 375.5330 0.0500 375.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 377.9330 1704.3000 378.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 377.9330 0.0500 378.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 382.7330 1704.3000 382.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 382.7330 0.0500 382.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 380.3330 1704.3000 380.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 380.3330 0.0500 380.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 387.5330 1704.3000 387.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 387.5330 0.0500 387.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 385.1330 1704.3000 385.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 385.1330 0.0500 385.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 389.9330 1704.3000 390.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 389.9330 0.0500 390.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 394.7330 1704.3000 394.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 394.7330 0.0500 394.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 392.3330 1704.3000 392.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 392.3330 0.0500 392.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 392.5060 1704.3000 399.5060 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 397.1330 1704.3000 397.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 397.1330 0.0500 397.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 399.5330 1704.3000 399.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 399.5330 0.0500 399.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 401.9330 1704.3000 402.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 401.9330 0.0500 402.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 404.3330 1704.3000 404.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 404.3330 0.0500 404.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 406.7330 1704.3000 406.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 406.7330 0.0500 406.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 409.1330 1704.3000 409.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 409.1330 0.0500 409.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 413.9330 1704.3000 414.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 413.9330 0.0500 414.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 411.5330 1704.3000 411.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 411.5330 0.0500 411.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 416.3330 1704.3000 416.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 416.3330 0.0500 416.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 418.7330 1704.3000 418.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 418.7330 0.0500 418.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 416.1340 1704.3000 423.1340 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 421.1330 1704.3000 421.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 421.1330 0.0500 421.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 423.5330 1704.3000 423.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 423.5330 0.0500 423.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 425.9330 1704.3000 426.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 425.9330 0.0500 426.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 428.3330 1704.3000 428.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 428.3330 0.0500 428.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 430.7330 1704.3000 430.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 430.7330 0.0500 430.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 433.1330 1704.3000 433.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 433.1330 0.0500 433.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 435.5330 1704.3000 435.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 435.5330 0.0500 435.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 437.9330 1704.3000 438.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 437.9330 0.0500 438.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 440.3330 1704.3000 440.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 440.3330 0.0500 440.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 442.7330 1704.3000 442.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 442.7330 0.0500 442.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 445.1330 1704.3000 445.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 445.1330 0.0500 445.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 439.7620 1704.3000 446.7620 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 447.5330 1704.3000 447.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 447.5330 0.0500 447.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 449.9330 1704.3000 450.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 449.9330 0.0500 450.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 452.3330 1704.3000 452.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 452.3330 0.0500 452.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 454.7330 1704.3000 454.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 454.7330 0.0500 454.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 457.1330 1704.3000 457.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 457.1330 0.0500 457.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 459.5330 1704.3000 459.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 459.5330 0.0500 459.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 461.9330 1704.3000 462.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 461.9330 0.0500 462.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 464.3330 1704.3000 464.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 464.3330 0.0500 464.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 463.3900 1704.3000 470.3900 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 469.1330 1704.3000 469.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 469.1330 0.0500 469.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 466.7330 1704.3000 466.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 466.7330 0.0500 466.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 471.5330 1704.3000 471.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 471.5330 0.0500 471.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 473.9330 1704.3000 474.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 473.9330 0.0500 474.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 476.3330 1704.3000 476.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 476.3330 0.0500 476.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 478.7330 1704.3000 478.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 478.7330 0.0500 478.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 481.1330 1704.3000 481.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 481.1330 0.0500 481.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 483.5330 1704.3000 483.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 483.5330 0.0500 483.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 485.9330 1704.3000 486.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 485.9330 0.0500 486.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 488.3330 1704.3000 488.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 488.3330 0.0500 488.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 487.0180 1704.3000 494.0180 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 490.7330 1704.3000 490.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 490.7330 0.0500 490.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 493.1330 1704.3000 493.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 493.1330 0.0500 493.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 495.5330 1704.3000 495.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 495.5330 0.0500 495.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 497.9330 1704.3000 498.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 497.9330 0.0500 498.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 500.3330 1704.3000 500.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 500.3330 0.0500 500.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 502.7330 1704.3000 502.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 502.7330 0.0500 502.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 505.1330 1704.3000 505.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 505.1330 0.0500 505.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 555.5330 1704.3000 555.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 555.5330 0.0500 555.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 560.3330 1704.3000 560.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 560.3330 0.0500 560.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 557.9330 1704.3000 558.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 557.9330 0.0500 558.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 558.8400 1704.3000 565.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 565.1330 1704.3000 565.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 565.1330 0.0500 565.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 562.7330 1704.3000 562.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 562.7330 0.0500 562.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 569.9330 1704.3000 570.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 569.9330 0.0500 570.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 567.5330 1704.3000 567.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 567.5330 0.0500 567.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 574.7330 1704.3000 574.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 574.7330 0.0500 574.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 572.3330 1704.3000 572.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 572.3330 0.0500 572.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 579.5330 1704.3000 579.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 579.5330 0.0500 579.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 577.1330 1704.3000 577.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 577.1330 0.0500 577.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 584.3330 1704.3000 584.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 584.3330 0.0500 584.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 581.9330 1704.3000 582.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 581.9330 0.0500 582.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 582.6540 1704.3000 589.6540 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 589.1330 1704.3000 589.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 589.1330 0.0500 589.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 586.7330 1704.3000 586.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 586.7330 0.0500 586.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 593.9330 1704.3000 594.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 593.9330 0.0500 594.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 591.5330 1704.3000 591.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 591.5330 0.0500 591.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 596.3330 1704.3000 596.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 596.3330 0.0500 596.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 601.1330 1704.3000 601.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 601.1330 0.0500 601.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 598.7330 1704.3000 598.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 598.7330 0.0500 598.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 605.9330 1704.3000 606.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 605.9330 0.0500 606.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 603.5330 1704.3000 603.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 603.5330 0.0500 603.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 606.2820 1704.3000 613.2820 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 610.7330 1704.3000 610.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 610.7330 0.0500 610.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 608.3330 1704.3000 608.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 608.3330 0.0500 608.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 615.5330 1704.3000 615.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 615.5330 0.0500 615.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 613.1330 1704.3000 613.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 613.1330 0.0500 613.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 617.9330 1704.3000 618.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 617.9330 0.0500 618.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 620.3330 1704.3000 620.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 620.3330 0.0500 620.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 625.1330 1704.3000 625.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 625.1330 0.0500 625.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 622.7330 1704.3000 622.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 622.7330 0.0500 622.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 629.9330 1704.3000 630.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 629.9330 0.0500 630.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 627.5330 1704.3000 627.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 627.5330 0.0500 627.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 634.7330 1704.3000 634.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 634.7330 0.0500 634.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 632.3330 1704.3000 632.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 632.3330 0.0500 632.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 629.9100 1704.3000 636.9100 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 637.1330 1704.3000 637.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 637.1330 0.0500 637.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 639.5330 1704.3000 639.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 639.5330 0.0500 639.6670 ;
    END
    PORT
      LAYER IA ;
        RECT 38.1210 0.0000 45.1210 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 38.1210 640.4000 45.1210 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 13.8110 0.0000 20.8110 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 13.8110 640.4000 20.8110 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 62.4310 0.0000 69.4310 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 62.4310 640.4000 69.4310 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 279.0550 0.0000 286.0550 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 279.0550 640.4000 286.0550 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 254.7450 0.0000 261.7450 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 254.7450 640.4000 261.7450 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 230.5900 0.0000 237.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 230.5900 640.4000 237.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 351.9850 0.0000 358.9850 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 351.9850 640.4000 358.9850 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 327.6750 0.0000 334.6750 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 327.6750 640.4000 334.6750 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 303.3650 0.0000 310.3650 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 303.3650 640.4000 310.3650 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 424.9150 0.0000 431.9150 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 424.9150 640.4000 431.9150 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 400.6050 0.0000 407.6050 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 400.6050 640.4000 407.6050 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 376.2950 0.0000 383.2950 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 376.2950 640.4000 383.2950 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 449.2250 0.0000 456.2250 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 449.2250 640.4000 456.2250 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 473.5350 0.0000 480.5350 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 473.5350 640.4000 480.5350 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 665.8490 0.0000 672.8490 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 665.8490 640.4000 672.8490 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 641.6940 0.0000 648.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 641.6940 640.4000 648.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 690.1590 0.0000 697.1590 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 690.1590 640.4000 697.1590 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 763.0890 0.0000 770.0890 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 763.0890 640.4000 770.0890 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 738.7790 0.0000 745.7790 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 738.7790 640.4000 745.7790 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 714.4690 0.0000 721.4690 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 714.4690 640.4000 721.4690 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 836.0190 0.0000 843.0190 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 836.0190 640.4000 843.0190 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 811.7090 0.0000 818.7090 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 811.7090 640.4000 818.7090 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 787.3990 0.0000 794.3990 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 787.3990 640.4000 794.3990 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 884.6390 0.0000 891.6390 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 884.6390 640.4000 891.6390 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 860.3290 0.0000 867.3290 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 860.3290 640.4000 867.3290 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1076.9530 0.0000 1083.9530 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1076.9530 640.4000 1083.9530 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1052.7980 0.0000 1059.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1052.7980 640.4000 1059.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1149.8830 0.0000 1156.8830 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1149.8830 640.4000 1156.8830 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1125.5730 0.0000 1132.5730 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1125.5730 640.4000 1132.5730 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1101.2630 0.0000 1108.2630 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1101.2630 640.4000 1108.2630 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1174.1930 0.0000 1181.1930 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1174.1930 640.4000 1181.1930 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1247.1230 0.0000 1254.1230 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1247.1230 640.4000 1254.1230 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1222.8130 0.0000 1229.8130 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1222.8130 640.4000 1229.8130 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1198.5030 0.0000 1205.5030 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1198.5030 640.4000 1205.5030 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1295.7430 0.0000 1302.7430 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1295.7430 640.4000 1302.7430 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1271.4330 0.0000 1278.4330 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1271.4330 640.4000 1278.4330 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1488.0570 0.0000 1495.0570 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1488.0570 640.4000 1495.0570 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1463.9020 0.0000 1470.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1463.9020 640.4000 1470.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1560.9870 0.0000 1567.9870 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1560.9870 640.4000 1567.9870 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1536.6770 0.0000 1543.6770 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1536.6770 640.4000 1543.6770 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1512.3670 0.0000 1519.3670 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1512.3670 640.4000 1519.3670 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1633.9170 0.0000 1640.9170 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1633.9170 640.4000 1640.9170 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1609.6070 0.0000 1616.6070 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1609.6070 640.4000 1616.6070 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1585.2970 0.0000 1592.2970 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1585.2970 640.4000 1592.2970 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 110.5900 0.0000 117.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 86.5900 0.0000 93.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 206.5900 0.0000 213.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 182.5900 0.0000 189.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 158.5900 0.0000 165.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 134.5900 0.0000 141.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 593.6940 0.0000 600.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 569.6940 0.0000 576.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 545.6940 0.0000 552.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 521.6940 0.0000 528.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 497.6940 0.0000 504.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 617.6940 0.0000 624.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1028.7980 0.0000 1035.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1004.7980 0.0000 1011.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 980.7980 0.0000 987.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 956.7980 0.0000 963.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 932.7980 0.0000 939.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 908.7980 0.0000 915.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1391.9020 0.0000 1398.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1367.9020 0.0000 1374.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1343.9020 0.0000 1350.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1319.9020 0.0000 1326.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1415.9020 0.0000 1422.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1439.9020 0.0000 1446.9020 0.4000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER LB ;
        RECT 1696.8600 136.2960 1704.3000 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 491.8400 1704.3000 521.8400 ;
    END
    PORT
      LAYER IA ;
        RECT 1427.9020 640.4000 1434.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1451.9020 640.4000 1458.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1331.9020 640.4000 1338.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1355.9020 640.4000 1362.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1379.9020 640.4000 1386.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1403.9020 640.4000 1410.9020 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 443.4480 1726.8600 521.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 554.3330 1704.3000 554.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 551.9330 1704.3000 552.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 549.5330 1704.3000 549.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 547.1330 1704.3000 547.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 544.7330 1704.3000 544.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 542.3330 1704.3000 542.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 539.9330 1704.3000 540.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 537.5330 1704.3000 537.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 535.1330 1704.3000 535.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 532.7330 1704.3000 532.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 530.3330 1704.3000 530.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 527.9330 1704.3000 528.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 1467.9020 546.8400 1704.3000 553.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1467.9020 522.8400 1704.3000 529.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 525.5330 1704.3000 525.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 523.1330 1704.3000 523.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 520.7330 1704.3000 520.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 518.3330 1704.3000 518.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 515.9330 1704.3000 516.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 513.5330 1704.3000 513.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 511.1330 1704.3000 511.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 508.7330 1704.3000 508.8670 ;
    END
    PORT
      LAYER LB ;
        RECT 1443.0160 428.4480 1506.3080 458.4480 ;
    END
    PORT
      LAYER LB ;
        RECT 1696.8600 87.9040 1726.8600 166.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 199.1330 1704.3000 199.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 196.7330 1704.3000 196.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 194.3330 1704.3000 194.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 191.9330 1704.3000 192.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 189.5330 1704.3000 189.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 187.1330 1704.3000 187.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 184.7330 1704.3000 184.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 1467.9020 191.2960 1704.3000 198.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 182.3330 1704.3000 182.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 179.9330 1704.3000 180.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 177.5330 1704.3000 177.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 175.1330 1704.3000 175.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 172.7330 1704.3000 172.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 170.3330 1704.3000 170.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 167.9330 1704.3000 168.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 165.5330 1704.3000 165.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 1467.9020 167.2960 1704.3000 174.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 163.1330 1704.3000 163.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 160.7330 1704.3000 160.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 158.3330 1704.3000 158.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 155.9330 1704.3000 156.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 153.5330 1704.3000 153.6670 ;
    END
    PORT
      LAYER LB ;
        RECT 1417.4020 454.0620 1447.4020 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1417.4020 98.5180 1447.4020 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1331.9020 491.8400 1361.9020 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 491.8400 1361.9020 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 443.4480 1315.7560 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1331.9020 136.2960 1361.9020 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 136.2960 1361.9020 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1285.7560 87.9040 1315.7560 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1443.0160 72.9040 1506.3080 102.9040 ;
    END
    PORT
      LAYER IB ;
        RECT 1056.7980 546.8400 1314.9020 553.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1056.7980 522.8400 1314.9020 529.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 1056.7980 191.2960 1314.9020 198.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 1056.7980 167.2960 1314.9020 174.2960 ;
    END
    PORT
      LAYER IA ;
        RECT 944.7980 640.4000 951.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 968.7980 640.4000 975.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 992.7980 640.4000 999.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1016.7980 640.4000 1023.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1040.7980 640.4000 1047.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 920.7980 640.4000 927.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 629.6940 640.4000 636.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 509.6940 640.4000 516.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 533.6940 640.4000 540.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 557.6940 640.4000 564.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 581.6940 640.4000 588.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 605.6940 640.4000 612.6940 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 1031.9120 428.4480 1095.2040 458.4480 ;
    END
    PORT
      LAYER LB ;
        RECT 1006.2980 454.0620 1036.2980 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 920.7980 491.8400 950.7980 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 491.8400 950.7980 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 443.4480 904.6520 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 1006.2980 98.5180 1036.2980 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 920.7980 136.2960 950.7980 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 136.2960 950.7980 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 874.6520 87.9040 904.6520 166.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 645.6940 546.8400 903.7980 553.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 645.6940 522.8400 903.7980 529.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 645.6940 191.2960 903.7980 198.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 645.6940 167.2960 903.7980 174.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 428.4480 625.1940 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 428.4480 670.1000 458.4480 ;
    END
    PORT
      LAYER LB ;
        RECT 509.6940 428.4480 539.6940 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 464.5470 428.4480 539.6940 458.4480 ;
    END
    PORT
      LAYER IB ;
        RECT 234.5900 546.8400 492.6940 553.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 234.5900 522.8400 492.6940 529.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 234.5900 191.2960 492.6940 198.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 234.5900 167.2960 492.6940 174.2960 ;
    END
    PORT
      LAYER IA ;
        RECT 146.5900 640.4000 153.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 170.5900 640.4000 177.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 194.5900 640.4000 201.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 218.5900 640.4000 225.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 98.5900 640.4000 105.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 122.5900 640.4000 129.5900 640.8000 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 428.4480 214.0900 521.8400 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 428.4480 258.9960 458.4480 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 554.3330 0.0500 554.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 551.9330 0.0500 552.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 549.5330 0.0500 549.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 547.1330 0.0500 547.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 544.7330 0.0500 544.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 542.3330 0.0500 542.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 539.9330 0.0500 540.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 537.5330 0.0500 537.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 535.1330 0.0500 535.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 532.7330 0.0500 532.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 530.3330 0.0500 530.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 527.9330 0.0500 528.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 525.5330 0.0500 525.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 523.1330 0.0500 523.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 520.7330 0.0500 520.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 518.3330 0.0500 518.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 515.9330 0.0500 516.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 513.5330 0.0500 513.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 511.1330 0.0500 511.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 508.7330 0.0500 508.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 522.8400 81.5900 529.8400 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 546.8400 81.5900 553.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 199.1330 0.0500 199.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 196.7330 0.0500 196.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 194.3330 0.0500 194.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 191.9330 0.0500 192.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 189.5330 0.0500 189.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 187.1330 0.0500 187.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 184.7330 0.0500 184.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 182.3330 0.0500 182.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 179.9330 0.0500 180.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 177.5330 0.0500 177.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 175.1330 0.0500 175.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 172.7330 0.0500 172.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 170.3330 0.0500 170.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 167.9330 0.0500 168.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 165.5330 0.0500 165.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 163.1330 0.0500 163.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 160.7330 0.0500 160.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 158.3330 0.0500 158.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 155.9330 0.0500 156.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 153.5330 0.0500 153.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 167.2960 81.5900 174.2960 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 191.2960 81.5900 198.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 1031.9120 72.9040 1095.2040 102.9040 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 72.9040 625.1940 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 595.1940 72.9040 670.1000 102.9040 ;
    END
    PORT
      LAYER LB ;
        RECT 509.6940 72.9040 539.6940 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 464.5470 72.9040 539.6940 102.9040 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 72.9040 214.0900 166.2960 ;
    END
    PORT
      LAYER LB ;
        RECT 184.0900 72.9040 258.9960 102.9040 ;
    END
    PORT
      LAYER IA ;
        RECT 1670.3820 0.0000 1677.3820 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1670.3820 640.4000 1677.3820 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1694.6920 0.0000 1701.6920 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1694.6920 640.4000 1701.6920 640.8000 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 -0.0670 1704.3000 0.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 1.5200 1704.3000 8.5200 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 2.3330 1704.3000 2.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 2.3330 0.0500 2.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 4.7330 1704.3000 4.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 4.7330 0.0500 4.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 7.1330 1704.3000 7.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 7.1330 0.0500 7.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 9.5330 1704.3000 9.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 9.5330 0.0500 9.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 11.9330 1704.3000 12.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 11.9330 0.0500 12.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 14.3330 1704.3000 14.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 14.3330 0.0500 14.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 16.7330 1704.3000 16.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 16.7330 0.0500 16.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 19.1330 1704.3000 19.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 19.1330 0.0500 19.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 21.5330 1704.3000 21.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 21.5330 0.0500 21.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 23.9330 1704.3000 24.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 23.9330 0.0500 24.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 26.3330 1704.3000 26.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 26.3330 0.0500 26.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 25.1480 1704.3000 32.1480 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 28.7330 1704.3000 28.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 28.7330 0.0500 28.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 31.1330 1704.3000 31.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 31.1330 0.0500 31.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 33.5330 1704.3000 33.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 33.5330 0.0500 33.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 35.9330 1704.3000 36.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 35.9330 0.0500 36.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 38.3330 1704.3000 38.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 38.3330 0.0500 38.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 40.7330 1704.3000 40.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 40.7330 0.0500 40.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 43.1330 1704.3000 43.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 43.1330 0.0500 43.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 45.5330 1704.3000 45.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 45.5330 0.0500 45.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 47.9330 1704.3000 48.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 47.9330 0.0500 48.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 50.3330 1704.3000 50.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 50.3330 0.0500 50.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 48.7760 1704.3000 55.7760 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 52.7330 1704.3000 52.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 52.7330 0.0500 52.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 55.1330 1704.3000 55.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 55.1330 0.0500 55.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 57.5330 1704.3000 57.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 57.5330 0.0500 57.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 59.9330 1704.3000 60.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 59.9330 0.0500 60.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 62.3330 1704.3000 62.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 62.3330 0.0500 62.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 64.7330 1704.3000 64.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 64.7330 0.0500 64.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 67.1330 1704.3000 67.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 67.1330 0.0500 67.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 69.5330 1704.3000 69.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 69.5330 0.0500 69.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 71.9330 1704.3000 72.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 71.9330 0.0500 72.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 72.4040 1704.3000 79.4040 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 74.3330 1704.3000 74.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 74.3330 0.0500 74.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 76.7330 1704.3000 76.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 76.7330 0.0500 76.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 79.1330 1704.3000 79.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 79.1330 0.0500 79.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 81.5330 1704.3000 81.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 81.5330 0.0500 81.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 83.9330 1704.3000 84.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 83.9330 0.0500 84.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 86.3330 1704.3000 86.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 86.3330 0.0500 86.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 88.7330 1704.3000 88.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 88.7330 0.0500 88.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 91.1330 1704.3000 91.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 91.1330 0.0500 91.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 93.5330 1704.3000 93.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 93.5330 0.0500 93.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 95.9330 1704.3000 96.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 95.9330 0.0500 96.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 96.0320 1704.3000 103.0320 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 98.3330 1704.3000 98.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 98.3330 0.0500 98.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 100.7330 1704.3000 100.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 100.7330 0.0500 100.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 103.1330 1704.3000 103.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 103.1330 0.0500 103.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 105.5330 1704.3000 105.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 105.5330 0.0500 105.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 107.9330 1704.3000 108.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 107.9330 0.0500 108.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 110.3330 1704.3000 110.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 110.3330 0.0500 110.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 112.7330 1704.3000 112.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 112.7330 0.0500 112.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 115.1330 1704.3000 115.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 115.1330 0.0500 115.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 117.5330 1704.3000 117.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 117.5330 0.0500 117.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 119.9330 1704.3000 120.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 119.9330 0.0500 120.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 122.3330 1704.3000 122.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 122.3330 0.0500 122.4670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 119.6600 1704.3000 126.6600 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 124.7330 1704.3000 124.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 124.7330 0.0500 124.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 127.1330 1704.3000 127.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 127.1330 0.0500 127.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 129.5330 1704.3000 129.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 129.5330 0.0500 129.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 131.9330 1704.3000 132.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 131.9330 0.0500 132.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 134.3330 1704.3000 134.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 134.3330 0.0500 134.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 136.7330 1704.3000 136.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 136.7330 0.0500 136.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 141.5330 1704.3000 141.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 141.5330 0.0500 141.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 139.1330 1704.3000 139.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 139.1330 0.0500 139.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 143.2960 1704.3000 150.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 143.9330 1704.3000 144.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 143.9330 0.0500 144.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 146.3330 1704.3000 146.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 146.3330 0.0500 146.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 151.1330 1704.3000 151.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 151.1330 0.0500 151.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 148.7330 1704.3000 148.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 148.7330 0.0500 148.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 201.5330 1704.3000 201.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 201.5330 0.0500 201.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 203.9330 1704.3000 204.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 203.9330 0.0500 204.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 206.3330 1704.3000 206.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 206.3330 0.0500 206.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 208.7330 1704.3000 208.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 208.7330 0.0500 208.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 213.5330 1704.3000 213.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 213.5330 0.0500 213.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 211.1330 1704.3000 211.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 211.1330 0.0500 211.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 218.3330 1704.3000 218.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 218.3330 0.0500 218.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 215.9330 1704.3000 216.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 215.9330 0.0500 216.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 215.2960 1704.3000 222.2960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 223.1330 1704.3000 223.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 223.1330 0.0500 223.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 220.7330 1704.3000 220.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 220.7330 0.0500 220.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 227.9330 1704.3000 228.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 227.9330 0.0500 228.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 225.5330 1704.3000 225.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 225.5330 0.0500 225.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 232.7330 1704.3000 232.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 232.7330 0.0500 232.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 230.3330 1704.3000 230.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 230.3330 0.0500 230.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 237.5330 1704.3000 237.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 237.5330 0.0500 237.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 235.1330 1704.3000 235.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 235.1330 0.0500 235.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 242.3330 1704.3000 242.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 242.3330 0.0500 242.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 239.9330 1704.3000 240.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 239.9330 0.0500 240.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 238.9240 1704.3000 245.9240 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 247.1330 1704.3000 247.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 247.1330 0.0500 247.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 244.7330 1704.3000 244.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 244.7330 0.0500 244.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 251.9330 1704.3000 252.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 251.9330 0.0500 252.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 249.5330 1704.3000 249.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 249.5330 0.0500 249.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 256.7330 1704.3000 256.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 256.7330 0.0500 256.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 254.3330 1704.3000 254.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 254.3330 0.0500 254.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 259.1330 1704.3000 259.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 259.1330 0.0500 259.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 263.9330 1704.3000 264.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 263.9330 0.0500 264.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 261.5330 1704.3000 261.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 261.5330 0.0500 261.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 262.5520 1704.3000 269.5520 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 268.7330 1704.3000 268.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 268.7330 0.0500 268.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 266.3330 1704.3000 266.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 266.3330 0.0500 266.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 273.5330 1704.3000 273.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 273.5330 0.0500 273.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 271.1330 1704.3000 271.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 271.1330 0.0500 271.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 278.3330 1704.3000 278.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 278.3330 0.0500 278.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 275.9330 1704.3000 276.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 275.9330 0.0500 276.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 283.1330 1704.3000 283.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 283.1330 0.0500 283.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 280.7330 1704.3000 280.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 280.7330 0.0500 280.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 287.9330 1704.3000 288.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 287.9330 0.0500 288.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 285.5330 1704.3000 285.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 285.5330 0.0500 285.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 286.1800 1704.3000 293.1800 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 292.7330 1704.3000 292.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 292.7330 0.0500 292.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 290.3330 1704.3000 290.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 290.3330 0.0500 290.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 297.5330 1704.3000 297.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 297.5330 0.0500 297.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 295.1330 1704.3000 295.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 295.1330 0.0500 295.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 302.3330 1704.3000 302.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 302.3330 0.0500 302.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 299.9330 1704.3000 300.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 299.9330 0.0500 300.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 307.1330 1704.3000 307.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 307.1330 0.0500 307.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 304.7330 1704.3000 304.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 304.7330 0.0500 304.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 314.3330 1704.3000 314.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 314.3330 0.0500 314.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 311.9330 1704.3000 312.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 311.9330 0.0500 312.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 309.5330 1704.3000 309.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 309.5330 0.0500 309.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 309.8080 1704.3000 316.8080 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 319.1330 1704.3000 319.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 319.1330 0.0500 319.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 316.7330 1704.3000 316.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 316.7330 0.0500 316.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 323.9330 1704.3000 324.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 323.9330 0.0500 324.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 321.5330 1704.3000 321.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 321.5330 0.0500 321.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 328.7330 1704.3000 328.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 328.7330 0.0500 328.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 326.3330 1704.3000 326.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 326.3330 0.0500 326.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 333.5330 1704.3000 333.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 333.5330 0.0500 333.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 331.1330 1704.3000 331.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 331.1330 0.0500 331.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 333.4360 1704.3000 340.4360 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 335.9330 1704.3000 336.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 335.9330 0.0500 336.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 338.3330 1704.3000 338.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 338.3330 0.0500 338.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 343.1330 1704.3000 343.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 343.1330 0.0500 343.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 340.7330 1704.3000 340.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 340.7330 0.0500 340.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 347.9330 1704.3000 348.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 347.9330 0.0500 348.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 345.5330 1704.3000 345.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 345.5330 0.0500 345.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 352.7330 1704.3000 352.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 352.7330 0.0500 352.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 350.3330 1704.3000 350.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 350.3330 0.0500 350.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 355.1330 1704.3000 355.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 355.1330 0.0500 355.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 357.5330 1704.3000 357.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 357.5330 0.0500 357.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 357.0640 1704.3000 364.0640 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 362.3330 1704.3000 362.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 362.3330 0.0500 362.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 359.9330 1704.3000 360.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 359.9330 0.0500 360.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 364.7330 1704.3000 364.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 364.7330 0.0500 364.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 369.5330 1704.3000 369.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 369.5330 0.0500 369.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 367.1330 1704.3000 367.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 367.1330 0.0500 367.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 374.3330 1704.3000 374.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 374.3330 0.0500 374.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 371.9330 1704.3000 372.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 371.9330 0.0500 372.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 379.1330 1704.3000 379.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 379.1330 0.0500 379.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 376.7330 1704.3000 376.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 376.7330 0.0500 376.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 383.9330 1704.3000 384.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 383.9330 0.0500 384.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 381.5330 1704.3000 381.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 381.5330 0.0500 381.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 380.6920 1704.3000 387.6920 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 388.7330 1704.3000 388.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 388.7330 0.0500 388.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 386.3330 1704.3000 386.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 386.3330 0.0500 386.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 393.5330 1704.3000 393.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 393.5330 0.0500 393.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 391.1330 1704.3000 391.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 391.1330 0.0500 391.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 398.3330 1704.3000 398.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 398.3330 0.0500 398.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 395.9330 1704.3000 396.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 395.9330 0.0500 396.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 403.1330 1704.3000 403.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 403.1330 0.0500 403.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 400.7330 1704.3000 400.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 400.7330 0.0500 400.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 404.3200 1704.3000 411.3200 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 407.9330 1704.3000 408.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 407.9330 0.0500 408.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 405.5330 1704.3000 405.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 405.5330 0.0500 405.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 412.7330 1704.3000 412.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 412.7330 0.0500 412.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 410.3330 1704.3000 410.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 410.3330 0.0500 410.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 415.1330 1704.3000 415.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 415.1330 0.0500 415.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 419.9330 1704.3000 420.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 419.9330 0.0500 420.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 417.5330 1704.3000 417.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 417.5330 0.0500 417.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 424.7330 1704.3000 424.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 424.7330 0.0500 424.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 422.3330 1704.3000 422.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 422.3330 0.0500 422.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 429.5330 1704.3000 429.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 429.5330 0.0500 429.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 427.1330 1704.3000 427.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 427.1330 0.0500 427.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 427.9480 1704.3000 434.9480 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 434.3330 1704.3000 434.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 434.3330 0.0500 434.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 431.9330 1704.3000 432.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 431.9330 0.0500 432.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 439.1330 1704.3000 439.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 439.1330 0.0500 439.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 436.7330 1704.3000 436.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 436.7330 0.0500 436.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 443.9330 1704.3000 444.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 443.9330 0.0500 444.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 441.5330 1704.3000 441.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 441.5330 0.0500 441.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 448.7330 1704.3000 448.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 448.7330 0.0500 448.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 446.3330 1704.3000 446.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 446.3330 0.0500 446.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 453.5330 1704.3000 453.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 453.5330 0.0500 453.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 451.1330 1704.3000 451.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 451.1330 0.0500 451.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 451.5760 1704.3000 458.5760 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 458.3330 1704.3000 458.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 458.3330 0.0500 458.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 455.9330 1704.3000 456.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 455.9330 0.0500 456.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 463.1330 1704.3000 463.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 463.1330 0.0500 463.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 460.7330 1704.3000 460.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 460.7330 0.0500 460.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 470.3330 1704.3000 470.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 470.3330 0.0500 470.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 467.9330 1704.3000 468.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 467.9330 0.0500 468.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 465.5330 1704.3000 465.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 465.5330 0.0500 465.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 472.7330 1704.3000 472.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 472.7330 0.0500 472.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 475.1330 1704.3000 475.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 475.1330 0.0500 475.2670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 475.2040 1704.3000 482.2040 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 477.5330 1704.3000 477.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 477.5330 0.0500 477.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 479.9330 1704.3000 480.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 479.9330 0.0500 480.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 482.3330 1704.3000 482.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 482.3330 0.0500 482.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 484.7330 1704.3000 484.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 484.7330 0.0500 484.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 487.1330 1704.3000 487.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 487.1330 0.0500 487.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 489.5330 1704.3000 489.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 489.5330 0.0500 489.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 491.9330 1704.3000 492.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 491.9330 0.0500 492.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 494.3330 1704.3000 494.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 494.3330 0.0500 494.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 496.7330 1704.3000 496.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 496.7330 0.0500 496.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 499.1330 1704.3000 499.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 499.1330 0.0500 499.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 501.5330 1704.3000 501.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 501.5330 0.0500 501.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 503.9330 1704.3000 504.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 503.9330 0.0500 504.0670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 498.8400 1704.3000 505.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 506.3330 1704.3000 506.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 506.3330 0.0500 506.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 559.1330 1704.3000 559.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 559.1330 0.0500 559.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 556.7330 1704.3000 556.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 556.7330 0.0500 556.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 563.9330 1704.3000 564.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 563.9330 0.0500 564.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 561.5330 1704.3000 561.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 561.5330 0.0500 561.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 568.7330 1704.3000 568.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 568.7330 0.0500 568.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 566.3330 1704.3000 566.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 566.3330 0.0500 566.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 571.1330 1704.3000 571.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 571.1330 0.0500 571.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 575.9330 1704.3000 576.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 575.9330 0.0500 576.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 573.5330 1704.3000 573.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 573.5330 0.0500 573.6670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 570.8400 1704.3000 577.8400 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 580.7330 1704.3000 580.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 580.7330 0.0500 580.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 578.3330 1704.3000 578.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 578.3330 0.0500 578.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 585.5330 1704.3000 585.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 585.5330 0.0500 585.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 583.1330 1704.3000 583.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 583.1330 0.0500 583.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 590.3330 1704.3000 590.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 590.3330 0.0500 590.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 587.9330 1704.3000 588.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 587.9330 0.0500 588.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 595.1330 1704.3000 595.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 595.1330 0.0500 595.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 592.7330 1704.3000 592.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 592.7330 0.0500 592.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 594.4680 1704.3000 601.4680 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 599.9330 1704.3000 600.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 599.9330 0.0500 600.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 597.5330 1704.3000 597.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 597.5330 0.0500 597.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 602.3330 1704.3000 602.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 602.3330 0.0500 602.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 604.7330 1704.3000 604.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 604.7330 0.0500 604.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 609.5330 1704.3000 609.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 609.5330 0.0500 609.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 607.1330 1704.3000 607.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 607.1330 0.0500 607.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 614.3330 1704.3000 614.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 614.3330 0.0500 614.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 611.9330 1704.3000 612.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 611.9330 0.0500 612.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 619.1330 1704.3000 619.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 619.1330 0.0500 619.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 616.7330 1704.3000 616.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 616.7330 0.0500 616.8670 ;
    END
    PORT
      LAYER IB ;
        RECT 0.0000 618.0960 1704.3000 625.0960 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 621.5330 1704.3000 621.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 621.5330 0.0500 621.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 626.3330 1704.3000 626.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 626.3330 0.0500 626.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 623.9330 1704.3000 624.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 623.9330 0.0500 624.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 631.1330 1704.3000 631.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 631.1330 0.0500 631.2670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 628.7330 1704.3000 628.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 628.7330 0.0500 628.8670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 635.9330 1704.3000 636.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 635.9330 0.0500 636.0670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 633.5330 1704.3000 633.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 633.5330 0.0500 633.6670 ;
    END
    PORT
      LAYER M2 ;
        RECT 1704.2500 638.3330 1704.3000 638.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 638.3330 0.0500 638.4670 ;
    END
    PORT
      LAYER M2 ;
        RECT 0.0000 640.7330 1704.3000 640.8670 ;
    END
    PORT
      LAYER IA ;
        RECT 1.6560 0.0000 8.6560 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1.6560 640.4000 8.6560 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 25.9660 0.0000 32.9660 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 25.9660 640.4000 32.9660 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 50.2760 0.0000 57.2760 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 50.2760 640.4000 57.2760 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 74.5900 0.0000 81.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 74.5900 640.4000 81.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 266.9000 0.0000 273.9000 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 266.9000 640.4000 273.9000 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 242.5900 0.0000 249.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 242.5900 640.4000 249.5900 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 364.1400 0.0000 371.1400 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 364.1400 640.4000 371.1400 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 339.8300 0.0000 346.8300 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 339.8300 640.4000 346.8300 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 315.5200 0.0000 322.5200 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 315.5200 640.4000 322.5200 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 291.2100 0.0000 298.2100 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 291.2100 640.4000 298.2100 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 437.0700 0.0000 444.0700 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 437.0700 640.4000 444.0700 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 412.7600 0.0000 419.7600 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 412.7600 640.4000 419.7600 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 388.4500 0.0000 395.4500 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 388.4500 640.4000 395.4500 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 461.3800 0.0000 468.3800 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 461.3800 640.4000 468.3800 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 485.6940 0.0000 492.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 485.6940 640.4000 492.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 678.0040 0.0000 685.0040 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 678.0040 640.4000 685.0040 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 653.6940 0.0000 660.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 653.6940 640.4000 660.6940 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 750.9340 0.0000 757.9340 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 750.9340 640.4000 757.9340 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 726.6240 0.0000 733.6240 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 726.6240 640.4000 733.6240 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 702.3140 0.0000 709.3140 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 702.3140 640.4000 709.3140 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 823.8640 0.0000 830.8640 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 823.8640 640.4000 830.8640 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 799.5540 0.0000 806.5540 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 799.5540 640.4000 806.5540 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 775.2440 0.0000 782.2440 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 775.2440 640.4000 782.2440 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 848.1740 0.0000 855.1740 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 848.1740 640.4000 855.1740 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 872.4840 0.0000 879.4840 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 872.4840 640.4000 879.4840 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 896.7980 0.0000 903.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 896.7980 640.4000 903.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1089.1080 0.0000 1096.1080 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1089.1080 640.4000 1096.1080 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1064.7980 0.0000 1071.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1064.7980 640.4000 1071.7980 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1162.0380 0.0000 1169.0380 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1162.0380 640.4000 1169.0380 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1137.7280 0.0000 1144.7280 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1137.7280 640.4000 1144.7280 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1113.4180 0.0000 1120.4180 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1113.4180 640.4000 1120.4180 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1234.9680 0.0000 1241.9680 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1234.9680 640.4000 1241.9680 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1210.6580 0.0000 1217.6580 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1210.6580 640.4000 1217.6580 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1186.3480 0.0000 1193.3480 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1186.3480 640.4000 1193.3480 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1283.5880 0.0000 1290.5880 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1283.5880 640.4000 1290.5880 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1259.2780 0.0000 1266.2780 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1259.2780 640.4000 1266.2780 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1307.9020 0.0000 1314.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1307.9020 640.4000 1314.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1475.9020 0.0000 1482.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1475.9020 640.4000 1482.9020 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1548.8320 0.0000 1555.8320 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1548.8320 640.4000 1555.8320 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1524.5220 0.0000 1531.5220 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1524.5220 640.4000 1531.5220 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1500.2120 0.0000 1507.2120 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1500.2120 640.4000 1507.2120 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1573.1420 0.0000 1580.1420 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1573.1420 640.4000 1580.1420 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1646.0720 0.0000 1653.0720 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1646.0720 640.4000 1653.0720 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1621.7620 0.0000 1628.7620 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1621.7620 640.4000 1628.7620 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 1597.4520 0.0000 1604.4520 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1597.4520 640.4000 1604.4520 640.8000 ;
    END
    PORT
      LAYER IA ;
        RECT 122.5900 0.0000 129.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 98.5900 0.0000 105.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 218.5900 0.0000 225.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 194.5900 0.0000 201.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 170.5900 0.0000 177.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 146.5900 0.0000 153.5900 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 605.6940 0.0000 612.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 581.6940 0.0000 588.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 557.6940 0.0000 564.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 533.6940 0.0000 540.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 509.6940 0.0000 516.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 629.6940 0.0000 636.6940 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1040.7980 0.0000 1047.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1016.7980 0.0000 1023.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 992.7980 0.0000 999.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 968.7980 0.0000 975.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 944.7980 0.0000 951.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 920.7980 0.0000 927.7980 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1403.9020 0.0000 1410.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1379.9020 0.0000 1386.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1355.9020 0.0000 1362.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1331.9020 0.0000 1338.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1451.9020 0.0000 1458.9020 0.4000 ;
    END
    PORT
      LAYER IA ;
        RECT 1427.9020 0.0000 1434.9020 0.4000 ;
    END
  END VDD
  OBS
    LAYER OVERLAP ;
    LAYER IB ;
      RECT 0.0000 0.0000 1704.3000 639.7240 ;
    LAYER IA ;
      RECT 0.0000 0.0000 3.0060 0.6000 ;
      RECT 7.3060 0.0000 27.3160 0.6000 ;
      RECT 31.6160 0.0000 51.6260 0.6000 ;
      RECT 55.9260 0.0000 75.9400 0.6000 ;
      RECT 80.2400 0.0000 99.9400 0.6000 ;
      RECT 104.2400 0.0000 123.9400 0.6000 ;
      RECT 128.2400 0.0000 147.9400 0.6000 ;
      RECT 152.2400 0.0000 171.9400 0.6000 ;
      RECT 176.2400 0.0000 195.9400 0.6000 ;
      RECT 200.2400 0.0000 219.9400 0.6000 ;
      RECT 224.2400 0.0000 243.9400 0.6000 ;
      RECT 248.2400 0.0000 268.2500 0.6000 ;
      RECT 272.5500 0.0000 292.5600 0.6000 ;
      RECT 296.8600 0.0000 316.8700 0.6000 ;
      RECT 321.1700 0.0000 341.1800 0.6000 ;
      RECT 345.4800 0.0000 365.4900 0.6000 ;
      RECT 369.7900 0.0000 389.8000 0.6000 ;
      RECT 394.1000 0.0000 414.1100 0.6000 ;
      RECT 418.4100 0.0000 438.4200 0.6000 ;
      RECT 442.7200 0.0000 462.7300 0.6000 ;
      RECT 467.0300 0.0000 487.0440 0.6000 ;
      RECT 491.3440 0.0000 511.0440 0.6000 ;
      RECT 515.3440 0.0000 535.0440 0.6000 ;
      RECT 539.3440 0.0000 559.0440 0.6000 ;
      RECT 563.3440 0.0000 583.0440 0.6000 ;
      RECT 587.3440 0.0000 607.0440 0.6000 ;
      RECT 611.3440 0.0000 631.0440 0.6000 ;
      RECT 635.3440 0.0000 655.0440 0.6000 ;
      RECT 659.3440 0.0000 679.3540 0.6000 ;
      RECT 683.6540 0.0000 703.6640 0.6000 ;
      RECT 707.9640 0.0000 727.9740 0.6000 ;
      RECT 732.2740 0.0000 752.2840 0.6000 ;
      RECT 756.5840 0.0000 776.5940 0.6000 ;
      RECT 780.8940 0.0000 800.9040 0.6000 ;
      RECT 805.2040 0.0000 825.2140 0.6000 ;
      RECT 829.5140 0.0000 849.5240 0.6000 ;
      RECT 853.8240 0.0000 873.8340 0.6000 ;
      RECT 878.1340 0.0000 898.1480 0.6000 ;
      RECT 902.4480 0.0000 922.1480 0.6000 ;
      RECT 926.4480 0.0000 946.1480 0.6000 ;
      RECT 950.4480 0.0000 970.1480 0.6000 ;
      RECT 974.4480 0.0000 994.1480 0.6000 ;
      RECT 998.4480 0.0000 1018.1480 0.6000 ;
      RECT 1022.4480 0.0000 1042.1480 0.6000 ;
      RECT 1046.4480 0.0000 1066.1480 0.6000 ;
      RECT 1070.4480 0.0000 1090.4580 0.6000 ;
      RECT 1094.7580 0.0000 1114.7680 0.6000 ;
      RECT 1119.0680 0.0000 1139.0780 0.6000 ;
      RECT 1143.3780 0.0000 1163.3880 0.6000 ;
      RECT 1167.6880 0.0000 1187.6980 0.6000 ;
      RECT 1191.9980 0.0000 1212.0080 0.6000 ;
      RECT 1216.3080 0.0000 1236.3180 0.6000 ;
      RECT 1240.6180 0.0000 1260.6280 0.6000 ;
      RECT 1264.9280 0.0000 1284.9380 0.6000 ;
      RECT 1289.2380 0.0000 1309.2520 0.6000 ;
      RECT 1313.5520 0.0000 1333.2520 0.6000 ;
      RECT 1337.5520 0.0000 1357.2520 0.6000 ;
      RECT 1361.5520 0.0000 1381.2520 0.6000 ;
      RECT 1385.5520 0.0000 1405.2520 0.6000 ;
      RECT 1409.5520 0.0000 1429.2520 0.6000 ;
      RECT 1433.5520 0.0000 1453.2520 0.6000 ;
      RECT 1457.5520 0.0000 1477.2520 0.6000 ;
      RECT 1481.5520 0.0000 1501.5620 0.6000 ;
      RECT 1505.8620 0.0000 1525.8720 0.6000 ;
      RECT 1530.1720 0.0000 1550.1820 0.6000 ;
      RECT 1554.4820 0.0000 1574.4920 0.6000 ;
      RECT 1578.7920 0.0000 1598.8020 0.6000 ;
      RECT 1603.1020 0.0000 1623.1120 0.6000 ;
      RECT 1627.4120 0.0000 1647.4220 0.6000 ;
      RECT 1651.7220 0.0000 1671.7320 0.6000 ;
      RECT 1676.0320 0.0000 1696.0420 0.6000 ;
      RECT 1700.3420 0.0000 1704.3000 0.6000 ;
      RECT 0.0000 0.6000 1704.3000 640.2000 ;
      RECT 0.0000 640.2000 3.0060 640.8000 ;
      RECT 7.3060 640.2000 27.3160 640.8000 ;
      RECT 31.6160 640.2000 51.6260 640.8000 ;
      RECT 55.9260 640.2000 75.9400 640.8000 ;
      RECT 80.2400 640.2000 99.9400 640.8000 ;
      RECT 104.2400 640.2000 123.9400 640.8000 ;
      RECT 128.2400 640.2000 147.9400 640.8000 ;
      RECT 152.2400 640.2000 171.9400 640.8000 ;
      RECT 176.2400 640.2000 195.9400 640.8000 ;
      RECT 200.2400 640.2000 219.9400 640.8000 ;
      RECT 224.2400 640.2000 243.9400 640.8000 ;
      RECT 248.2400 640.2000 268.2500 640.8000 ;
      RECT 272.5500 640.2000 292.5600 640.8000 ;
      RECT 296.8600 640.2000 316.8700 640.8000 ;
      RECT 321.1700 640.2000 341.1800 640.8000 ;
      RECT 345.4800 640.2000 365.4900 640.8000 ;
      RECT 369.7900 640.2000 389.8000 640.8000 ;
      RECT 394.1000 640.2000 414.1100 640.8000 ;
      RECT 418.4100 640.2000 438.4200 640.8000 ;
      RECT 442.7200 640.2000 462.7300 640.8000 ;
      RECT 467.0300 640.2000 487.0440 640.8000 ;
      RECT 491.3440 640.2000 511.0440 640.8000 ;
      RECT 515.3440 640.2000 535.0440 640.8000 ;
      RECT 539.3440 640.2000 559.0440 640.8000 ;
      RECT 563.3440 640.2000 583.0440 640.8000 ;
      RECT 587.3440 640.2000 607.0440 640.8000 ;
      RECT 611.3440 640.2000 631.0440 640.8000 ;
      RECT 635.3440 640.2000 655.0440 640.8000 ;
      RECT 659.3440 640.2000 679.3540 640.8000 ;
      RECT 683.6540 640.2000 703.6640 640.8000 ;
      RECT 707.9640 640.2000 727.9740 640.8000 ;
      RECT 732.2740 640.2000 752.2840 640.8000 ;
      RECT 756.5840 640.2000 776.5940 640.8000 ;
      RECT 780.8940 640.2000 800.9040 640.8000 ;
      RECT 805.2040 640.2000 825.2140 640.8000 ;
      RECT 829.5140 640.2000 849.5240 640.8000 ;
      RECT 853.8240 640.2000 873.8340 640.8000 ;
      RECT 878.1340 640.2000 898.1480 640.8000 ;
      RECT 902.4480 640.2000 922.1480 640.8000 ;
      RECT 926.4480 640.2000 946.1480 640.8000 ;
      RECT 950.4480 640.2000 970.1480 640.8000 ;
      RECT 974.4480 640.2000 994.1480 640.8000 ;
      RECT 998.4480 640.2000 1018.1480 640.8000 ;
      RECT 1022.4480 640.2000 1042.1480 640.8000 ;
      RECT 1046.4480 640.2000 1066.1480 640.8000 ;
      RECT 1070.4480 640.2000 1090.4580 640.8000 ;
      RECT 1094.7580 640.2000 1114.7680 640.8000 ;
      RECT 1119.0680 640.2000 1139.0780 640.8000 ;
      RECT 1143.3780 640.2000 1163.3880 640.8000 ;
      RECT 1167.6880 640.2000 1187.6980 640.8000 ;
      RECT 1191.9980 640.2000 1212.0080 640.8000 ;
      RECT 1216.3080 640.2000 1236.3180 640.8000 ;
      RECT 1240.6180 640.2000 1260.6280 640.8000 ;
      RECT 1264.9280 640.2000 1284.9380 640.8000 ;
      RECT 1289.2380 640.2000 1309.2520 640.8000 ;
      RECT 1313.5520 640.2000 1333.2520 640.8000 ;
      RECT 1337.5520 640.2000 1357.2520 640.8000 ;
      RECT 1361.5520 640.2000 1381.2520 640.8000 ;
      RECT 1385.5520 640.2000 1405.2520 640.8000 ;
      RECT 1409.5520 640.2000 1429.2520 640.8000 ;
      RECT 1433.5520 640.2000 1453.2520 640.8000 ;
      RECT 1457.5520 640.2000 1477.2520 640.8000 ;
      RECT 1481.5520 640.2000 1501.5620 640.8000 ;
      RECT 1505.8620 640.2000 1525.8720 640.8000 ;
      RECT 1530.1720 640.2000 1550.1820 640.8000 ;
      RECT 1554.4820 640.2000 1574.4920 640.8000 ;
      RECT 1578.7920 640.2000 1598.8020 640.8000 ;
      RECT 1603.1020 640.2000 1623.1120 640.8000 ;
      RECT 1627.4120 640.2000 1647.4220 640.8000 ;
      RECT 1651.7220 640.2000 1671.7320 640.8000 ;
      RECT 1676.0320 640.2000 1696.0420 640.8000 ;
      RECT 1700.3420 640.2000 1704.3000 640.8000 ;
    LAYER B2 ;
      RECT 0.0000 0.0000 3.3060 0.1670 ;
      RECT 7.0060 0.0000 27.6160 0.1670 ;
      RECT 31.3160 0.0000 51.9260 0.1670 ;
      RECT 55.6260 0.0000 76.2400 0.1670 ;
      RECT 79.9400 0.0000 100.2400 0.1670 ;
      RECT 103.9400 0.0000 124.2400 0.1670 ;
      RECT 127.9400 0.0000 148.2400 0.1670 ;
      RECT 151.9400 0.0000 172.2400 0.1670 ;
      RECT 175.9400 0.0000 196.2400 0.1670 ;
      RECT 199.9400 0.0000 220.2400 0.1670 ;
      RECT 223.9400 0.0000 244.2400 0.1670 ;
      RECT 247.9400 0.0000 268.5500 0.1670 ;
      RECT 272.2500 0.0000 292.8600 0.1670 ;
      RECT 296.5600 0.0000 317.1700 0.1670 ;
      RECT 320.8700 0.0000 341.4800 0.1670 ;
      RECT 345.1800 0.0000 365.7900 0.1670 ;
      RECT 369.4900 0.0000 390.1000 0.1670 ;
      RECT 393.8000 0.0000 414.4100 0.1670 ;
      RECT 418.1100 0.0000 438.7200 0.1670 ;
      RECT 442.4200 0.0000 463.0300 0.1670 ;
      RECT 466.7300 0.0000 487.3440 0.1670 ;
      RECT 491.0440 0.0000 511.3440 0.1670 ;
      RECT 515.0440 0.0000 535.3440 0.1670 ;
      RECT 539.0440 0.0000 559.3440 0.1670 ;
      RECT 563.0440 0.0000 583.3440 0.1670 ;
      RECT 587.0440 0.0000 607.3440 0.1670 ;
      RECT 611.0440 0.0000 631.3440 0.1670 ;
      RECT 635.0440 0.0000 655.3440 0.1670 ;
      RECT 659.0440 0.0000 679.6540 0.1670 ;
      RECT 683.3540 0.0000 703.9640 0.1670 ;
      RECT 707.6640 0.0000 728.2740 0.1670 ;
      RECT 731.9740 0.0000 752.5840 0.1670 ;
      RECT 756.2840 0.0000 776.8940 0.1670 ;
      RECT 780.5940 0.0000 801.2040 0.1670 ;
      RECT 804.9040 0.0000 825.5140 0.1670 ;
      RECT 829.2140 0.0000 849.8240 0.1670 ;
      RECT 853.5240 0.0000 874.1340 0.1670 ;
      RECT 877.8340 0.0000 898.4480 0.1670 ;
      RECT 902.1480 0.0000 922.4480 0.1670 ;
      RECT 926.1480 0.0000 946.4480 0.1670 ;
      RECT 950.1480 0.0000 970.4480 0.1670 ;
      RECT 974.1480 0.0000 994.4480 0.1670 ;
      RECT 998.1480 0.0000 1018.4480 0.1670 ;
      RECT 1022.1480 0.0000 1042.4480 0.1670 ;
      RECT 1046.1480 0.0000 1066.4480 0.1670 ;
      RECT 1070.1480 0.0000 1090.7580 0.1670 ;
      RECT 1094.4580 0.0000 1115.0680 0.1670 ;
      RECT 1118.7680 0.0000 1139.3780 0.1670 ;
      RECT 1143.0780 0.0000 1163.6880 0.1670 ;
      RECT 1167.3880 0.0000 1187.9980 0.1670 ;
      RECT 1191.6980 0.0000 1212.3080 0.1670 ;
      RECT 1216.0080 0.0000 1236.6180 0.1670 ;
      RECT 1240.3180 0.0000 1260.9280 0.1670 ;
      RECT 1264.6280 0.0000 1285.2380 0.1670 ;
      RECT 1288.9380 0.0000 1309.5520 0.1670 ;
      RECT 1313.2520 0.0000 1333.5520 0.1670 ;
      RECT 1337.2520 0.0000 1357.5520 0.1670 ;
      RECT 1361.2520 0.0000 1381.5520 0.1670 ;
      RECT 1385.2520 0.0000 1405.5520 0.1670 ;
      RECT 1409.2520 0.0000 1429.5520 0.1670 ;
      RECT 1433.2520 0.0000 1453.5520 0.1670 ;
      RECT 1457.2520 0.0000 1477.5520 0.1670 ;
      RECT 1481.2520 0.0000 1501.8620 0.1670 ;
      RECT 1505.5620 0.0000 1526.1720 0.1670 ;
      RECT 1529.8720 0.0000 1550.4820 0.1670 ;
      RECT 1554.1820 0.0000 1574.7920 0.1670 ;
      RECT 1578.4920 0.0000 1599.1020 0.1670 ;
      RECT 1602.8020 0.0000 1623.4120 0.1670 ;
      RECT 1627.1120 0.0000 1647.7220 0.1670 ;
      RECT 1651.4220 0.0000 1672.0320 0.1670 ;
      RECT 1675.7320 0.0000 1696.3420 0.1670 ;
      RECT 0.0000 0.1670 3.3060 0.3000 ;
      RECT 7.0060 0.1670 27.6160 0.3000 ;
      RECT 31.3160 0.1670 51.9260 0.3000 ;
      RECT 55.6260 0.1670 76.2400 0.3000 ;
      RECT 79.9400 0.1670 100.2400 0.3000 ;
      RECT 103.9400 0.1670 124.2400 0.3000 ;
      RECT 127.9400 0.1670 148.2400 0.3000 ;
      RECT 151.9400 0.1670 172.2400 0.3000 ;
      RECT 175.9400 0.1670 196.2400 0.3000 ;
      RECT 199.9400 0.1670 220.2400 0.3000 ;
      RECT 223.9400 0.1670 244.2400 0.3000 ;
      RECT 247.9400 0.1670 268.5500 0.3000 ;
      RECT 272.2500 0.1670 292.8600 0.3000 ;
      RECT 296.5600 0.1670 317.1700 0.3000 ;
      RECT 320.8700 0.1670 341.4800 0.3000 ;
      RECT 345.1800 0.1670 365.7900 0.3000 ;
      RECT 369.4900 0.1670 390.1000 0.3000 ;
      RECT 393.8000 0.1670 414.4100 0.3000 ;
      RECT 418.1100 0.1670 438.7200 0.3000 ;
      RECT 442.4200 0.1670 463.0300 0.3000 ;
      RECT 466.7300 0.1670 487.3440 0.3000 ;
      RECT 491.0440 0.1670 511.3440 0.3000 ;
      RECT 515.0440 0.1670 535.3440 0.3000 ;
      RECT 539.0440 0.1670 559.3440 0.3000 ;
      RECT 563.0440 0.1670 583.3440 0.3000 ;
      RECT 587.0440 0.1670 607.3440 0.3000 ;
      RECT 611.0440 0.1670 631.3440 0.3000 ;
      RECT 635.0440 0.1670 655.3440 0.3000 ;
      RECT 659.0440 0.1670 679.6540 0.3000 ;
      RECT 683.3540 0.1670 703.9640 0.3000 ;
      RECT 707.6640 0.1670 728.2740 0.3000 ;
      RECT 731.9740 0.1670 752.5840 0.3000 ;
      RECT 756.2840 0.1670 776.8940 0.3000 ;
      RECT 780.5940 0.1670 801.2040 0.3000 ;
      RECT 804.9040 0.1670 825.5140 0.3000 ;
      RECT 829.2140 0.1670 849.8240 0.3000 ;
      RECT 853.5240 0.1670 874.1340 0.3000 ;
      RECT 877.8340 0.1670 898.4480 0.3000 ;
      RECT 902.1480 0.1670 922.4480 0.3000 ;
      RECT 926.1480 0.1670 946.4480 0.3000 ;
      RECT 950.1480 0.1670 970.4480 0.3000 ;
      RECT 974.1480 0.1670 994.4480 0.3000 ;
      RECT 998.1480 0.1670 1018.4480 0.3000 ;
      RECT 1022.1480 0.1670 1042.4480 0.3000 ;
      RECT 1046.1480 0.1670 1066.4480 0.3000 ;
      RECT 1070.1480 0.1670 1090.7580 0.3000 ;
      RECT 1094.4580 0.1670 1115.0680 0.3000 ;
      RECT 1118.7680 0.1670 1139.3780 0.3000 ;
      RECT 1143.0780 0.1670 1163.6880 0.3000 ;
      RECT 1167.3880 0.1670 1187.9980 0.3000 ;
      RECT 1191.6980 0.1670 1212.3080 0.3000 ;
      RECT 1216.0080 0.1670 1236.6180 0.3000 ;
      RECT 1240.3180 0.1670 1260.9280 0.3000 ;
      RECT 1264.6280 0.1670 1285.2380 0.3000 ;
      RECT 1288.9380 0.1670 1309.5520 0.3000 ;
      RECT 1313.2520 0.1670 1333.5520 0.3000 ;
      RECT 1337.2520 0.1670 1357.5520 0.3000 ;
      RECT 1361.2520 0.1670 1381.5520 0.3000 ;
      RECT 1385.2520 0.1670 1405.5520 0.3000 ;
      RECT 1409.2520 0.1670 1429.5520 0.3000 ;
      RECT 1433.2520 0.1670 1453.5520 0.3000 ;
      RECT 1457.2520 0.1670 1477.5520 0.3000 ;
      RECT 1481.2520 0.1670 1501.8620 0.3000 ;
      RECT 1505.5620 0.1670 1526.1720 0.3000 ;
      RECT 1529.8720 0.1670 1550.4820 0.3000 ;
      RECT 1554.1820 0.1670 1574.7920 0.3000 ;
      RECT 1578.4920 0.1670 1599.1020 0.3000 ;
      RECT 1602.8020 0.1670 1623.4120 0.3000 ;
      RECT 1627.1120 0.1670 1647.7220 0.3000 ;
      RECT 1651.4220 0.1670 1672.0320 0.3000 ;
      RECT 1675.7320 0.1670 1696.3420 0.3000 ;
      RECT 1700.0420 0.0000 1704.3000 0.3000 ;
      RECT 0.0000 0.3000 1704.3000 640.5000 ;
      RECT 7.0060 640.5000 27.6160 640.6330 ;
      RECT 31.3160 640.5000 51.9260 640.6330 ;
      RECT 55.6260 640.5000 76.2400 640.6330 ;
      RECT 79.9400 640.5000 100.2400 640.6330 ;
      RECT 103.9400 640.5000 124.2400 640.6330 ;
      RECT 127.9400 640.5000 148.2400 640.6330 ;
      RECT 151.9400 640.5000 172.2400 640.6330 ;
      RECT 175.9400 640.5000 196.2400 640.6330 ;
      RECT 199.9400 640.5000 220.2400 640.6330 ;
      RECT 223.9400 640.5000 244.2400 640.6330 ;
      RECT 247.9400 640.5000 268.5500 640.6330 ;
      RECT 272.2500 640.5000 292.8600 640.6330 ;
      RECT 296.5600 640.5000 317.1700 640.6330 ;
      RECT 320.8700 640.5000 341.4800 640.6330 ;
      RECT 345.1800 640.5000 365.7900 640.6330 ;
      RECT 369.4900 640.5000 390.1000 640.6330 ;
      RECT 393.8000 640.5000 414.4100 640.6330 ;
      RECT 418.1100 640.5000 438.7200 640.6330 ;
      RECT 442.4200 640.5000 463.0300 640.6330 ;
      RECT 466.7300 640.5000 487.3440 640.6330 ;
      RECT 491.0440 640.5000 511.3440 640.6330 ;
      RECT 515.0440 640.5000 535.3440 640.6330 ;
      RECT 539.0440 640.5000 559.3440 640.6330 ;
      RECT 563.0440 640.5000 583.3440 640.6330 ;
      RECT 587.0440 640.5000 607.3440 640.6330 ;
      RECT 611.0440 640.5000 631.3440 640.6330 ;
      RECT 635.0440 640.5000 655.3440 640.6330 ;
      RECT 659.0440 640.5000 679.6540 640.6330 ;
      RECT 683.3540 640.5000 703.9640 640.6330 ;
      RECT 707.6640 640.5000 728.2740 640.6330 ;
      RECT 731.9740 640.5000 752.5840 640.6330 ;
      RECT 756.2840 640.5000 776.8940 640.6330 ;
      RECT 780.5940 640.5000 801.2040 640.6330 ;
      RECT 804.9040 640.5000 825.5140 640.6330 ;
      RECT 829.2140 640.5000 849.8240 640.6330 ;
      RECT 853.5240 640.5000 874.1340 640.6330 ;
      RECT 877.8340 640.5000 898.4480 640.6330 ;
      RECT 902.1480 640.5000 922.4480 640.6330 ;
      RECT 926.1480 640.5000 946.4480 640.6330 ;
      RECT 950.1480 640.5000 970.4480 640.6330 ;
      RECT 974.1480 640.5000 994.4480 640.6330 ;
      RECT 998.1480 640.5000 1018.4480 640.6330 ;
      RECT 1022.1480 640.5000 1042.4480 640.6330 ;
      RECT 1046.1480 640.5000 1066.4480 640.6330 ;
      RECT 1070.1480 640.5000 1090.7580 640.6330 ;
      RECT 1094.4580 640.5000 1115.0680 640.6330 ;
      RECT 1118.7680 640.5000 1139.3780 640.6330 ;
      RECT 1143.0780 640.5000 1163.6880 640.6330 ;
      RECT 1167.3880 640.5000 1187.9980 640.6330 ;
      RECT 1191.6980 640.5000 1212.3080 640.6330 ;
      RECT 1216.0080 640.5000 1236.6180 640.6330 ;
      RECT 1240.3180 640.5000 1260.9280 640.6330 ;
      RECT 1264.6280 640.5000 1285.2380 640.6330 ;
      RECT 1288.9380 640.5000 1309.5520 640.6330 ;
      RECT 1313.2520 640.5000 1333.5520 640.6330 ;
      RECT 1337.2520 640.5000 1357.5520 640.6330 ;
      RECT 1361.2520 640.5000 1381.5520 640.6330 ;
      RECT 1385.2520 640.5000 1405.5520 640.6330 ;
      RECT 1409.2520 640.5000 1429.5520 640.6330 ;
      RECT 1433.2520 640.5000 1453.5520 640.6330 ;
      RECT 1457.2520 640.5000 1477.5520 640.6330 ;
      RECT 1481.2520 640.5000 1501.8620 640.6330 ;
      RECT 1505.5620 640.5000 1526.1720 640.6330 ;
      RECT 1529.8720 640.5000 1550.4820 640.6330 ;
      RECT 1554.1820 640.5000 1574.7920 640.6330 ;
      RECT 1578.4920 640.5000 1599.1020 640.6330 ;
      RECT 1602.8020 640.5000 1623.4120 640.6330 ;
      RECT 1627.1120 640.5000 1647.7220 640.6330 ;
      RECT 1651.4220 640.5000 1672.0320 640.6330 ;
      RECT 1675.7320 640.5000 1696.3420 640.6330 ;
      RECT 1700.0420 640.5000 1704.3000 640.6330 ;
      RECT 0.0000 640.5000 3.3060 640.8000 ;
      RECT 7.0060 640.6330 27.6160 640.8000 ;
      RECT 31.3160 640.6330 51.9260 640.8000 ;
      RECT 55.6260 640.6330 76.2400 640.8000 ;
      RECT 79.9400 640.6330 100.2400 640.8000 ;
      RECT 103.9400 640.6330 124.2400 640.8000 ;
      RECT 127.9400 640.6330 148.2400 640.8000 ;
      RECT 151.9400 640.6330 172.2400 640.8000 ;
      RECT 175.9400 640.6330 196.2400 640.8000 ;
      RECT 199.9400 640.6330 220.2400 640.8000 ;
      RECT 223.9400 640.6330 244.2400 640.8000 ;
      RECT 247.9400 640.6330 268.5500 640.8000 ;
      RECT 272.2500 640.6330 292.8600 640.8000 ;
      RECT 296.5600 640.6330 317.1700 640.8000 ;
      RECT 320.8700 640.6330 341.4800 640.8000 ;
      RECT 345.1800 640.6330 365.7900 640.8000 ;
      RECT 369.4900 640.6330 390.1000 640.8000 ;
      RECT 393.8000 640.6330 414.4100 640.8000 ;
      RECT 418.1100 640.6330 438.7200 640.8000 ;
      RECT 442.4200 640.6330 463.0300 640.8000 ;
      RECT 466.7300 640.6330 487.3440 640.8000 ;
      RECT 491.0440 640.6330 511.3440 640.8000 ;
      RECT 515.0440 640.6330 535.3440 640.8000 ;
      RECT 539.0440 640.6330 559.3440 640.8000 ;
      RECT 563.0440 640.6330 583.3440 640.8000 ;
      RECT 587.0440 640.6330 607.3440 640.8000 ;
      RECT 611.0440 640.6330 631.3440 640.8000 ;
      RECT 635.0440 640.6330 655.3440 640.8000 ;
      RECT 659.0440 640.6330 679.6540 640.8000 ;
      RECT 683.3540 640.6330 703.9640 640.8000 ;
      RECT 707.6640 640.6330 728.2740 640.8000 ;
      RECT 731.9740 640.6330 752.5840 640.8000 ;
      RECT 756.2840 640.6330 776.8940 640.8000 ;
      RECT 780.5940 640.6330 801.2040 640.8000 ;
      RECT 804.9040 640.6330 825.5140 640.8000 ;
      RECT 829.2140 640.6330 849.8240 640.8000 ;
      RECT 853.5240 640.6330 874.1340 640.8000 ;
      RECT 877.8340 640.6330 898.4480 640.8000 ;
      RECT 902.1480 640.6330 922.4480 640.8000 ;
      RECT 926.1480 640.6330 946.4480 640.8000 ;
      RECT 950.1480 640.6330 970.4480 640.8000 ;
      RECT 974.1480 640.6330 994.4480 640.8000 ;
      RECT 998.1480 640.6330 1018.4480 640.8000 ;
      RECT 1022.1480 640.6330 1042.4480 640.8000 ;
      RECT 1046.1480 640.6330 1066.4480 640.8000 ;
      RECT 1070.1480 640.6330 1090.7580 640.8000 ;
      RECT 1094.4580 640.6330 1115.0680 640.8000 ;
      RECT 1118.7680 640.6330 1139.3780 640.8000 ;
      RECT 1143.0780 640.6330 1163.6880 640.8000 ;
      RECT 1167.3880 640.6330 1187.9980 640.8000 ;
      RECT 1191.6980 640.6330 1212.3080 640.8000 ;
      RECT 1216.0080 640.6330 1236.6180 640.8000 ;
      RECT 1240.3180 640.6330 1260.9280 640.8000 ;
      RECT 1264.6280 640.6330 1285.2380 640.8000 ;
      RECT 1288.9380 640.6330 1309.5520 640.8000 ;
      RECT 1313.2520 640.6330 1333.5520 640.8000 ;
      RECT 1337.2520 640.6330 1357.5520 640.8000 ;
      RECT 1361.2520 640.6330 1381.5520 640.8000 ;
      RECT 1385.2520 640.6330 1405.5520 640.8000 ;
      RECT 1409.2520 640.6330 1429.5520 640.8000 ;
      RECT 1433.2520 640.6330 1453.5520 640.8000 ;
      RECT 1457.2520 640.6330 1477.5520 640.8000 ;
      RECT 1481.2520 640.6330 1501.8620 640.8000 ;
      RECT 1505.5620 640.6330 1526.1720 640.8000 ;
      RECT 1529.8720 640.6330 1550.4820 640.8000 ;
      RECT 1554.1820 640.6330 1574.7920 640.8000 ;
      RECT 1578.4920 640.6330 1599.1020 640.8000 ;
      RECT 1602.8020 640.6330 1623.4120 640.8000 ;
      RECT 1627.1120 640.6330 1647.7220 640.8000 ;
      RECT 1651.4220 640.6330 1672.0320 640.8000 ;
      RECT 1675.7320 640.6330 1696.3420 640.8000 ;
      RECT 1700.0420 640.6330 1704.3000 640.8000 ;
    LAYER B1 ;
      RECT 7.0060 0.0000 27.6160 0.1670 ;
      RECT 0.0000 0.0000 3.3060 0.1670 ;
      RECT 31.3160 0.0000 51.9260 0.1670 ;
      RECT 55.6260 0.0000 76.2400 0.1670 ;
      RECT 79.9400 0.0000 100.2400 0.1670 ;
      RECT 103.9400 0.0000 124.2400 0.1670 ;
      RECT 127.9400 0.0000 148.2400 0.1670 ;
      RECT 151.9400 0.0000 172.2400 0.1670 ;
      RECT 175.9400 0.0000 196.2400 0.1670 ;
      RECT 199.9400 0.0000 220.2400 0.1670 ;
      RECT 223.9400 0.0000 244.2400 0.1670 ;
      RECT 247.9400 0.0000 268.5500 0.1670 ;
      RECT 272.2500 0.0000 292.8600 0.1670 ;
      RECT 296.5600 0.0000 317.1700 0.1670 ;
      RECT 320.8700 0.0000 341.4800 0.1670 ;
      RECT 345.1800 0.0000 365.7900 0.1670 ;
      RECT 369.4900 0.0000 390.1000 0.1670 ;
      RECT 393.8000 0.0000 414.4100 0.1670 ;
      RECT 418.1100 0.0000 438.7200 0.1670 ;
      RECT 442.4200 0.0000 463.0300 0.1670 ;
      RECT 466.7300 0.0000 487.3440 0.1670 ;
      RECT 491.0440 0.0000 511.3440 0.1670 ;
      RECT 515.0440 0.0000 535.3440 0.1670 ;
      RECT 539.0440 0.0000 559.3440 0.1670 ;
      RECT 563.0440 0.0000 583.3440 0.1670 ;
      RECT 587.0440 0.0000 607.3440 0.1670 ;
      RECT 611.0440 0.0000 631.3440 0.1670 ;
      RECT 635.0440 0.0000 655.3440 0.1670 ;
      RECT 659.0440 0.0000 679.6540 0.1670 ;
      RECT 683.3540 0.0000 703.9640 0.1670 ;
      RECT 707.6640 0.0000 728.2740 0.1670 ;
      RECT 731.9740 0.0000 752.5840 0.1670 ;
      RECT 756.2840 0.0000 776.8940 0.1670 ;
      RECT 780.5940 0.0000 801.2040 0.1670 ;
      RECT 804.9040 0.0000 825.5140 0.1670 ;
      RECT 829.2140 0.0000 849.8240 0.1670 ;
      RECT 853.5240 0.0000 874.1340 0.1670 ;
      RECT 877.8340 0.0000 898.4480 0.1670 ;
      RECT 902.1480 0.0000 922.4480 0.1670 ;
      RECT 926.1480 0.0000 946.4480 0.1670 ;
      RECT 950.1480 0.0000 970.4480 0.1670 ;
      RECT 974.1480 0.0000 994.4480 0.1670 ;
      RECT 998.1480 0.0000 1018.4480 0.1670 ;
      RECT 1022.1480 0.0000 1042.4480 0.1670 ;
      RECT 1046.1480 0.0000 1066.4480 0.1670 ;
      RECT 1070.1480 0.0000 1090.7580 0.1670 ;
      RECT 1094.4580 0.0000 1115.0680 0.1670 ;
      RECT 1118.7680 0.0000 1139.3780 0.1670 ;
      RECT 1143.0780 0.0000 1163.6880 0.1670 ;
      RECT 1167.3880 0.0000 1187.9980 0.1670 ;
      RECT 1191.6980 0.0000 1212.3080 0.1670 ;
      RECT 1216.0080 0.0000 1236.6180 0.1670 ;
      RECT 1240.3180 0.0000 1260.9280 0.1670 ;
      RECT 1264.6280 0.0000 1285.2380 0.1670 ;
      RECT 1288.9380 0.0000 1309.5520 0.1670 ;
      RECT 1313.2520 0.0000 1333.5520 0.1670 ;
      RECT 1337.2520 0.0000 1357.5520 0.1670 ;
      RECT 1361.2520 0.0000 1381.5520 0.1670 ;
      RECT 1385.2520 0.0000 1405.5520 0.1670 ;
      RECT 1409.2520 0.0000 1429.5520 0.1670 ;
      RECT 1433.2520 0.0000 1453.5520 0.1670 ;
      RECT 1457.2520 0.0000 1477.5520 0.1670 ;
      RECT 1481.2520 0.0000 1501.8620 0.1670 ;
      RECT 1505.5620 0.0000 1526.1720 0.1670 ;
      RECT 1529.8720 0.0000 1550.4820 0.1670 ;
      RECT 1554.1820 0.0000 1574.7920 0.1670 ;
      RECT 1578.4920 0.0000 1599.1020 0.1670 ;
      RECT 1602.8020 0.0000 1623.4120 0.1670 ;
      RECT 1627.1120 0.0000 1647.7220 0.1670 ;
      RECT 1651.4220 0.0000 1672.0320 0.1670 ;
      RECT 1675.7320 0.0000 1696.3420 0.1670 ;
      RECT 1700.0420 0.0000 1704.3000 0.1670 ;
      RECT 0.0000 0.1670 1704.3000 640.6330 ;
      RECT 7.0060 640.6330 27.6160 640.8000 ;
      RECT 0.0000 640.6330 3.3060 640.8000 ;
      RECT 31.3160 640.6330 51.9260 640.8000 ;
      RECT 55.6260 640.6330 76.2400 640.8000 ;
      RECT 79.9400 640.6330 100.2400 640.8000 ;
      RECT 103.9400 640.6330 124.2400 640.8000 ;
      RECT 127.9400 640.6330 148.2400 640.8000 ;
      RECT 151.9400 640.6330 172.2400 640.8000 ;
      RECT 175.9400 640.6330 196.2400 640.8000 ;
      RECT 199.9400 640.6330 220.2400 640.8000 ;
      RECT 223.9400 640.6330 244.2400 640.8000 ;
      RECT 247.9400 640.6330 268.5500 640.8000 ;
      RECT 272.2500 640.6330 292.8600 640.8000 ;
      RECT 296.5600 640.6330 317.1700 640.8000 ;
      RECT 320.8700 640.6330 341.4800 640.8000 ;
      RECT 345.1800 640.6330 365.7900 640.8000 ;
      RECT 369.4900 640.6330 390.1000 640.8000 ;
      RECT 393.8000 640.6330 414.4100 640.8000 ;
      RECT 418.1100 640.6330 438.7200 640.8000 ;
      RECT 442.4200 640.6330 463.0300 640.8000 ;
      RECT 466.7300 640.6330 487.3440 640.8000 ;
      RECT 491.0440 640.6330 511.3440 640.8000 ;
      RECT 515.0440 640.6330 535.3440 640.8000 ;
      RECT 539.0440 640.6330 559.3440 640.8000 ;
      RECT 563.0440 640.6330 583.3440 640.8000 ;
      RECT 587.0440 640.6330 607.3440 640.8000 ;
      RECT 611.0440 640.6330 631.3440 640.8000 ;
      RECT 635.0440 640.6330 655.3440 640.8000 ;
      RECT 659.0440 640.6330 679.6540 640.8000 ;
      RECT 683.3540 640.6330 703.9640 640.8000 ;
      RECT 707.6640 640.6330 728.2740 640.8000 ;
      RECT 731.9740 640.6330 752.5840 640.8000 ;
      RECT 756.2840 640.6330 776.8940 640.8000 ;
      RECT 780.5940 640.6330 801.2040 640.8000 ;
      RECT 804.9040 640.6330 825.5140 640.8000 ;
      RECT 829.2140 640.6330 849.8240 640.8000 ;
      RECT 853.5240 640.6330 874.1340 640.8000 ;
      RECT 877.8340 640.6330 898.4480 640.8000 ;
      RECT 902.1480 640.6330 922.4480 640.8000 ;
      RECT 926.1480 640.6330 946.4480 640.8000 ;
      RECT 950.1480 640.6330 970.4480 640.8000 ;
      RECT 974.1480 640.6330 994.4480 640.8000 ;
      RECT 998.1480 640.6330 1018.4480 640.8000 ;
      RECT 1022.1480 640.6330 1042.4480 640.8000 ;
      RECT 1046.1480 640.6330 1066.4480 640.8000 ;
      RECT 1070.1480 640.6330 1090.7580 640.8000 ;
      RECT 1094.4580 640.6330 1115.0680 640.8000 ;
      RECT 1118.7680 640.6330 1139.3780 640.8000 ;
      RECT 1143.0780 640.6330 1163.6880 640.8000 ;
      RECT 1167.3880 640.6330 1187.9980 640.8000 ;
      RECT 1191.6980 640.6330 1212.3080 640.8000 ;
      RECT 1216.0080 640.6330 1236.6180 640.8000 ;
      RECT 1240.3180 640.6330 1260.9280 640.8000 ;
      RECT 1264.6280 640.6330 1285.2380 640.8000 ;
      RECT 1288.9380 640.6330 1309.5520 640.8000 ;
      RECT 1313.2520 640.6330 1333.5520 640.8000 ;
      RECT 1337.2520 640.6330 1357.5520 640.8000 ;
      RECT 1361.2520 640.6330 1381.5520 640.8000 ;
      RECT 1385.2520 640.6330 1405.5520 640.8000 ;
      RECT 1409.2520 640.6330 1429.5520 640.8000 ;
      RECT 1433.2520 640.6330 1453.5520 640.8000 ;
      RECT 1457.2520 640.6330 1477.5520 640.8000 ;
      RECT 1481.2520 640.6330 1501.8620 640.8000 ;
      RECT 1505.5620 640.6330 1526.1720 640.8000 ;
      RECT 1529.8720 640.6330 1550.4820 640.8000 ;
      RECT 1554.1820 640.6330 1574.7920 640.8000 ;
      RECT 1578.4920 640.6330 1599.1020 640.8000 ;
      RECT 1602.8020 640.6330 1623.4120 640.8000 ;
      RECT 1627.1120 640.6330 1647.7220 640.8000 ;
      RECT 1651.4220 640.6330 1672.0320 640.8000 ;
      RECT 1675.7320 640.6330 1696.3420 640.8000 ;
      RECT 1700.0420 640.6330 1704.3000 640.8000 ;
    LAYER M6 ;
      RECT 6.9560 0.0000 27.6660 0.1170 ;
      RECT 0.0000 0.0000 3.3560 0.1170 ;
      RECT 31.2660 0.0000 51.9760 0.1170 ;
      RECT 55.5760 0.0000 76.2900 0.1170 ;
      RECT 79.8900 0.0000 100.2900 0.1170 ;
      RECT 103.8900 0.0000 124.2900 0.1170 ;
      RECT 127.8900 0.0000 148.2900 0.1170 ;
      RECT 151.8900 0.0000 172.2900 0.1170 ;
      RECT 175.8900 0.0000 196.2900 0.1170 ;
      RECT 199.8900 0.0000 220.2900 0.1170 ;
      RECT 223.8900 0.0000 244.2900 0.1170 ;
      RECT 247.8900 0.0000 268.6000 0.1170 ;
      RECT 272.2000 0.0000 292.9100 0.1170 ;
      RECT 296.5100 0.0000 317.2200 0.1170 ;
      RECT 320.8200 0.0000 341.5300 0.1170 ;
      RECT 345.1300 0.0000 365.8400 0.1170 ;
      RECT 369.4400 0.0000 390.1500 0.1170 ;
      RECT 393.7500 0.0000 414.4600 0.1170 ;
      RECT 418.0600 0.0000 438.7700 0.1170 ;
      RECT 442.3700 0.0000 463.0800 0.1170 ;
      RECT 466.6800 0.0000 487.3940 0.1170 ;
      RECT 490.9940 0.0000 511.3940 0.1170 ;
      RECT 514.9940 0.0000 535.3940 0.1170 ;
      RECT 538.9940 0.0000 559.3940 0.1170 ;
      RECT 562.9940 0.0000 583.3940 0.1170 ;
      RECT 586.9940 0.0000 607.3940 0.1170 ;
      RECT 610.9940 0.0000 631.3940 0.1170 ;
      RECT 634.9940 0.0000 655.3940 0.1170 ;
      RECT 658.9940 0.0000 679.7040 0.1170 ;
      RECT 683.3040 0.0000 704.0140 0.1170 ;
      RECT 707.6140 0.0000 728.3240 0.1170 ;
      RECT 731.9240 0.0000 752.6340 0.1170 ;
      RECT 756.2340 0.0000 776.9440 0.1170 ;
      RECT 780.5440 0.0000 801.2540 0.1170 ;
      RECT 804.8540 0.0000 825.5640 0.1170 ;
      RECT 829.1640 0.0000 849.8740 0.1170 ;
      RECT 853.4740 0.0000 874.1840 0.1170 ;
      RECT 877.7840 0.0000 898.4980 0.1170 ;
      RECT 902.0980 0.0000 922.4980 0.1170 ;
      RECT 926.0980 0.0000 946.4980 0.1170 ;
      RECT 950.0980 0.0000 970.4980 0.1170 ;
      RECT 974.0980 0.0000 994.4980 0.1170 ;
      RECT 998.0980 0.0000 1018.4980 0.1170 ;
      RECT 1022.0980 0.0000 1042.4980 0.1170 ;
      RECT 1046.0980 0.0000 1066.4980 0.1170 ;
      RECT 1070.0980 0.0000 1090.8080 0.1170 ;
      RECT 1094.4080 0.0000 1115.1180 0.1170 ;
      RECT 1118.7180 0.0000 1139.4280 0.1170 ;
      RECT 1143.0280 0.0000 1163.7380 0.1170 ;
      RECT 1167.3380 0.0000 1188.0480 0.1170 ;
      RECT 1191.6480 0.0000 1212.3580 0.1170 ;
      RECT 1215.9580 0.0000 1236.6680 0.1170 ;
      RECT 1240.2680 0.0000 1260.9780 0.1170 ;
      RECT 1264.5780 0.0000 1285.2880 0.1170 ;
      RECT 1288.8880 0.0000 1309.6020 0.1170 ;
      RECT 1313.2020 0.0000 1333.6020 0.1170 ;
      RECT 1337.2020 0.0000 1357.6020 0.1170 ;
      RECT 1361.2020 0.0000 1381.6020 0.1170 ;
      RECT 1385.2020 0.0000 1405.6020 0.1170 ;
      RECT 1409.2020 0.0000 1429.6020 0.1170 ;
      RECT 1433.2020 0.0000 1453.6020 0.1170 ;
      RECT 1457.2020 0.0000 1477.6020 0.1170 ;
      RECT 1481.2020 0.0000 1501.9120 0.1170 ;
      RECT 1505.5120 0.0000 1526.2220 0.1170 ;
      RECT 1529.8220 0.0000 1550.5320 0.1170 ;
      RECT 1554.1320 0.0000 1574.8420 0.1170 ;
      RECT 1578.4420 0.0000 1599.1520 0.1170 ;
      RECT 1602.7520 0.0000 1623.4620 0.1170 ;
      RECT 1627.0620 0.0000 1647.7720 0.1170 ;
      RECT 1651.3720 0.0000 1672.0820 0.1170 ;
      RECT 1675.6820 0.0000 1696.3920 0.1170 ;
      RECT 1699.9920 0.0000 1704.3000 0.1170 ;
      RECT 0.0000 0.1170 1704.3000 640.6830 ;
      RECT 6.9560 640.6830 27.6660 640.8000 ;
      RECT 0.0000 640.6830 3.3560 640.8000 ;
      RECT 31.2660 640.6830 51.9760 640.8000 ;
      RECT 55.5760 640.6830 76.2900 640.8000 ;
      RECT 79.8900 640.6830 100.2900 640.8000 ;
      RECT 103.8900 640.6830 124.2900 640.8000 ;
      RECT 127.8900 640.6830 148.2900 640.8000 ;
      RECT 151.8900 640.6830 172.2900 640.8000 ;
      RECT 175.8900 640.6830 196.2900 640.8000 ;
      RECT 199.8900 640.6830 220.2900 640.8000 ;
      RECT 223.8900 640.6830 244.2900 640.8000 ;
      RECT 247.8900 640.6830 268.6000 640.8000 ;
      RECT 272.2000 640.6830 292.9100 640.8000 ;
      RECT 296.5100 640.6830 317.2200 640.8000 ;
      RECT 320.8200 640.6830 341.5300 640.8000 ;
      RECT 345.1300 640.6830 365.8400 640.8000 ;
      RECT 369.4400 640.6830 390.1500 640.8000 ;
      RECT 393.7500 640.6830 414.4600 640.8000 ;
      RECT 418.0600 640.6830 438.7700 640.8000 ;
      RECT 442.3700 640.6830 463.0800 640.8000 ;
      RECT 466.6800 640.6830 487.3940 640.8000 ;
      RECT 490.9940 640.6830 511.3940 640.8000 ;
      RECT 514.9940 640.6830 535.3940 640.8000 ;
      RECT 538.9940 640.6830 559.3940 640.8000 ;
      RECT 562.9940 640.6830 583.3940 640.8000 ;
      RECT 586.9940 640.6830 607.3940 640.8000 ;
      RECT 610.9940 640.6830 631.3940 640.8000 ;
      RECT 634.9940 640.6830 655.3940 640.8000 ;
      RECT 658.9940 640.6830 679.7040 640.8000 ;
      RECT 683.3040 640.6830 704.0140 640.8000 ;
      RECT 707.6140 640.6830 728.3240 640.8000 ;
      RECT 731.9240 640.6830 752.6340 640.8000 ;
      RECT 756.2340 640.6830 776.9440 640.8000 ;
      RECT 780.5440 640.6830 801.2540 640.8000 ;
      RECT 804.8540 640.6830 825.5640 640.8000 ;
      RECT 829.1640 640.6830 849.8740 640.8000 ;
      RECT 853.4740 640.6830 874.1840 640.8000 ;
      RECT 877.7840 640.6830 898.4980 640.8000 ;
      RECT 902.0980 640.6830 922.4980 640.8000 ;
      RECT 926.0980 640.6830 946.4980 640.8000 ;
      RECT 950.0980 640.6830 970.4980 640.8000 ;
      RECT 974.0980 640.6830 994.4980 640.8000 ;
      RECT 998.0980 640.6830 1018.4980 640.8000 ;
      RECT 1022.0980 640.6830 1042.4980 640.8000 ;
      RECT 1046.0980 640.6830 1066.4980 640.8000 ;
      RECT 1070.0980 640.6830 1090.8080 640.8000 ;
      RECT 1094.4080 640.6830 1115.1180 640.8000 ;
      RECT 1118.7180 640.6830 1139.4280 640.8000 ;
      RECT 1143.0280 640.6830 1163.7380 640.8000 ;
      RECT 1167.3380 640.6830 1188.0480 640.8000 ;
      RECT 1191.6480 640.6830 1212.3580 640.8000 ;
      RECT 1215.9580 640.6830 1236.6680 640.8000 ;
      RECT 1240.2680 640.6830 1260.9780 640.8000 ;
      RECT 1264.5780 640.6830 1285.2880 640.8000 ;
      RECT 1288.8880 640.6830 1309.6020 640.8000 ;
      RECT 1313.2020 640.6830 1333.6020 640.8000 ;
      RECT 1337.2020 640.6830 1357.6020 640.8000 ;
      RECT 1361.2020 640.6830 1381.6020 640.8000 ;
      RECT 1385.2020 640.6830 1405.6020 640.8000 ;
      RECT 1409.2020 640.6830 1429.6020 640.8000 ;
      RECT 1433.2020 640.6830 1453.6020 640.8000 ;
      RECT 1457.2020 640.6830 1477.6020 640.8000 ;
      RECT 1481.2020 640.6830 1501.9120 640.8000 ;
      RECT 1505.5120 640.6830 1526.2220 640.8000 ;
      RECT 1529.8220 640.6830 1550.5320 640.8000 ;
      RECT 1554.1320 640.6830 1574.8420 640.8000 ;
      RECT 1578.4420 640.6830 1599.1520 640.8000 ;
      RECT 1602.7520 640.6830 1623.4620 640.8000 ;
      RECT 1627.0620 640.6830 1647.7720 640.8000 ;
      RECT 1651.3720 640.6830 1672.0820 640.8000 ;
      RECT 1675.6820 640.6830 1696.3920 640.8000 ;
      RECT 1699.9920 640.6830 1704.3000 640.8000 ;
    LAYER M5 ;
      RECT 6.9560 0.0000 27.6660 0.1170 ;
      RECT 0.0000 0.0000 3.3560 0.1170 ;
      RECT 31.2660 0.0000 51.9760 0.1170 ;
      RECT 55.5760 0.0000 76.2900 0.1170 ;
      RECT 79.8900 0.0000 100.2900 0.1170 ;
      RECT 103.8900 0.0000 124.2900 0.1170 ;
      RECT 127.8900 0.0000 148.2900 0.1170 ;
      RECT 151.8900 0.0000 172.2900 0.1170 ;
      RECT 175.8900 0.0000 196.2900 0.1170 ;
      RECT 199.8900 0.0000 220.2900 0.1170 ;
      RECT 223.8900 0.0000 244.2900 0.1170 ;
      RECT 247.8900 0.0000 268.6000 0.1170 ;
      RECT 272.2000 0.0000 292.9100 0.1170 ;
      RECT 296.5100 0.0000 317.2200 0.1170 ;
      RECT 320.8200 0.0000 341.5300 0.1170 ;
      RECT 345.1300 0.0000 365.8400 0.1170 ;
      RECT 369.4400 0.0000 390.1500 0.1170 ;
      RECT 393.7500 0.0000 414.4600 0.1170 ;
      RECT 418.0600 0.0000 438.7700 0.1170 ;
      RECT 442.3700 0.0000 463.0800 0.1170 ;
      RECT 466.6800 0.0000 487.3940 0.1170 ;
      RECT 490.9940 0.0000 511.3940 0.1170 ;
      RECT 514.9940 0.0000 535.3940 0.1170 ;
      RECT 538.9940 0.0000 559.3940 0.1170 ;
      RECT 562.9940 0.0000 583.3940 0.1170 ;
      RECT 586.9940 0.0000 607.3940 0.1170 ;
      RECT 610.9940 0.0000 631.3940 0.1170 ;
      RECT 634.9940 0.0000 655.3940 0.1170 ;
      RECT 658.9940 0.0000 679.7040 0.1170 ;
      RECT 683.3040 0.0000 704.0140 0.1170 ;
      RECT 707.6140 0.0000 728.3240 0.1170 ;
      RECT 731.9240 0.0000 752.6340 0.1170 ;
      RECT 756.2340 0.0000 776.9440 0.1170 ;
      RECT 780.5440 0.0000 801.2540 0.1170 ;
      RECT 804.8540 0.0000 825.5640 0.1170 ;
      RECT 829.1640 0.0000 849.8740 0.1170 ;
      RECT 853.4740 0.0000 874.1840 0.1170 ;
      RECT 877.7840 0.0000 898.4980 0.1170 ;
      RECT 902.0980 0.0000 922.4980 0.1170 ;
      RECT 926.0980 0.0000 946.4980 0.1170 ;
      RECT 950.0980 0.0000 970.4980 0.1170 ;
      RECT 974.0980 0.0000 994.4980 0.1170 ;
      RECT 998.0980 0.0000 1018.4980 0.1170 ;
      RECT 1022.0980 0.0000 1042.4980 0.1170 ;
      RECT 1046.0980 0.0000 1066.4980 0.1170 ;
      RECT 1070.0980 0.0000 1090.8080 0.1170 ;
      RECT 1094.4080 0.0000 1115.1180 0.1170 ;
      RECT 1118.7180 0.0000 1139.4280 0.1170 ;
      RECT 1143.0280 0.0000 1163.7380 0.1170 ;
      RECT 1167.3380 0.0000 1188.0480 0.1170 ;
      RECT 1191.6480 0.0000 1212.3580 0.1170 ;
      RECT 1215.9580 0.0000 1236.6680 0.1170 ;
      RECT 1240.2680 0.0000 1260.9780 0.1170 ;
      RECT 1264.5780 0.0000 1285.2880 0.1170 ;
      RECT 1288.8880 0.0000 1309.6020 0.1170 ;
      RECT 1313.2020 0.0000 1333.6020 0.1170 ;
      RECT 1337.2020 0.0000 1357.6020 0.1170 ;
      RECT 1361.2020 0.0000 1381.6020 0.1170 ;
      RECT 1385.2020 0.0000 1405.6020 0.1170 ;
      RECT 1409.2020 0.0000 1429.6020 0.1170 ;
      RECT 1433.2020 0.0000 1453.6020 0.1170 ;
      RECT 1457.2020 0.0000 1477.6020 0.1170 ;
      RECT 1481.2020 0.0000 1501.9120 0.1170 ;
      RECT 1505.5120 0.0000 1526.2220 0.1170 ;
      RECT 1529.8220 0.0000 1550.5320 0.1170 ;
      RECT 1554.1320 0.0000 1574.8420 0.1170 ;
      RECT 1578.4420 0.0000 1599.1520 0.1170 ;
      RECT 1602.7520 0.0000 1623.4620 0.1170 ;
      RECT 1627.0620 0.0000 1647.7720 0.1170 ;
      RECT 1651.3720 0.0000 1672.0820 0.1170 ;
      RECT 1675.6820 0.0000 1696.3920 0.1170 ;
      RECT 1699.9920 0.0000 1704.3000 0.1170 ;
      RECT 0.0000 0.1170 1704.3000 640.6830 ;
      RECT 6.9560 640.6830 27.6660 640.8000 ;
      RECT 0.0000 640.6830 3.3560 640.8000 ;
      RECT 31.2660 640.6830 51.9760 640.8000 ;
      RECT 55.5760 640.6830 76.2900 640.8000 ;
      RECT 79.8900 640.6830 100.2900 640.8000 ;
      RECT 103.8900 640.6830 124.2900 640.8000 ;
      RECT 127.8900 640.6830 148.2900 640.8000 ;
      RECT 151.8900 640.6830 172.2900 640.8000 ;
      RECT 175.8900 640.6830 196.2900 640.8000 ;
      RECT 199.8900 640.6830 220.2900 640.8000 ;
      RECT 223.8900 640.6830 244.2900 640.8000 ;
      RECT 247.8900 640.6830 268.6000 640.8000 ;
      RECT 272.2000 640.6830 292.9100 640.8000 ;
      RECT 296.5100 640.6830 317.2200 640.8000 ;
      RECT 320.8200 640.6830 341.5300 640.8000 ;
      RECT 345.1300 640.6830 365.8400 640.8000 ;
      RECT 369.4400 640.6830 390.1500 640.8000 ;
      RECT 393.7500 640.6830 414.4600 640.8000 ;
      RECT 418.0600 640.6830 438.7700 640.8000 ;
      RECT 442.3700 640.6830 463.0800 640.8000 ;
      RECT 466.6800 640.6830 487.3940 640.8000 ;
      RECT 490.9940 640.6830 511.3940 640.8000 ;
      RECT 514.9940 640.6830 535.3940 640.8000 ;
      RECT 538.9940 640.6830 559.3940 640.8000 ;
      RECT 562.9940 640.6830 583.3940 640.8000 ;
      RECT 586.9940 640.6830 607.3940 640.8000 ;
      RECT 610.9940 640.6830 631.3940 640.8000 ;
      RECT 634.9940 640.6830 655.3940 640.8000 ;
      RECT 658.9940 640.6830 679.7040 640.8000 ;
      RECT 683.3040 640.6830 704.0140 640.8000 ;
      RECT 707.6140 640.6830 728.3240 640.8000 ;
      RECT 731.9240 640.6830 752.6340 640.8000 ;
      RECT 756.2340 640.6830 776.9440 640.8000 ;
      RECT 780.5440 640.6830 801.2540 640.8000 ;
      RECT 804.8540 640.6830 825.5640 640.8000 ;
      RECT 829.1640 640.6830 849.8740 640.8000 ;
      RECT 853.4740 640.6830 874.1840 640.8000 ;
      RECT 877.7840 640.6830 898.4980 640.8000 ;
      RECT 902.0980 640.6830 922.4980 640.8000 ;
      RECT 926.0980 640.6830 946.4980 640.8000 ;
      RECT 950.0980 640.6830 970.4980 640.8000 ;
      RECT 974.0980 640.6830 994.4980 640.8000 ;
      RECT 998.0980 640.6830 1018.4980 640.8000 ;
      RECT 1022.0980 640.6830 1042.4980 640.8000 ;
      RECT 1046.0980 640.6830 1066.4980 640.8000 ;
      RECT 1070.0980 640.6830 1090.8080 640.8000 ;
      RECT 1094.4080 640.6830 1115.1180 640.8000 ;
      RECT 1118.7180 640.6830 1139.4280 640.8000 ;
      RECT 1143.0280 640.6830 1163.7380 640.8000 ;
      RECT 1167.3380 640.6830 1188.0480 640.8000 ;
      RECT 1191.6480 640.6830 1212.3580 640.8000 ;
      RECT 1215.9580 640.6830 1236.6680 640.8000 ;
      RECT 1240.2680 640.6830 1260.9780 640.8000 ;
      RECT 1264.5780 640.6830 1285.2880 640.8000 ;
      RECT 1288.8880 640.6830 1309.6020 640.8000 ;
      RECT 1313.2020 640.6830 1333.6020 640.8000 ;
      RECT 1337.2020 640.6830 1357.6020 640.8000 ;
      RECT 1361.2020 640.6830 1381.6020 640.8000 ;
      RECT 1385.2020 640.6830 1405.6020 640.8000 ;
      RECT 1409.2020 640.6830 1429.6020 640.8000 ;
      RECT 1433.2020 640.6830 1453.6020 640.8000 ;
      RECT 1457.2020 640.6830 1477.6020 640.8000 ;
      RECT 1481.2020 640.6830 1501.9120 640.8000 ;
      RECT 1505.5120 640.6830 1526.2220 640.8000 ;
      RECT 1529.8220 640.6830 1550.5320 640.8000 ;
      RECT 1554.1320 640.6830 1574.8420 640.8000 ;
      RECT 1578.4420 640.6830 1599.1520 640.8000 ;
      RECT 1602.7520 640.6830 1623.4620 640.8000 ;
      RECT 1627.0620 640.6830 1647.7720 640.8000 ;
      RECT 1651.3720 640.6830 1672.0820 640.8000 ;
      RECT 1675.6820 640.6830 1696.3920 640.8000 ;
      RECT 1699.9920 640.6830 1704.3000 640.8000 ;
    LAYER M4 ;
      RECT 6.9560 0.0000 27.6660 0.1170 ;
      RECT 0.0000 0.0000 3.3560 0.1170 ;
      RECT 31.2660 0.0000 51.9760 0.1170 ;
      RECT 55.5760 0.0000 76.2900 0.1170 ;
      RECT 79.8900 0.0000 100.2900 0.1170 ;
      RECT 103.8900 0.0000 124.2900 0.1170 ;
      RECT 127.8900 0.0000 148.2900 0.1170 ;
      RECT 151.8900 0.0000 172.2900 0.1170 ;
      RECT 175.8900 0.0000 196.2900 0.1170 ;
      RECT 199.8900 0.0000 220.2900 0.1170 ;
      RECT 223.8900 0.0000 244.2900 0.1170 ;
      RECT 247.8900 0.0000 268.6000 0.1170 ;
      RECT 272.2000 0.0000 292.9100 0.1170 ;
      RECT 296.5100 0.0000 317.2200 0.1170 ;
      RECT 320.8200 0.0000 341.5300 0.1170 ;
      RECT 345.1300 0.0000 365.8400 0.1170 ;
      RECT 369.4400 0.0000 390.1500 0.1170 ;
      RECT 393.7500 0.0000 414.4600 0.1170 ;
      RECT 418.0600 0.0000 438.7700 0.1170 ;
      RECT 442.3700 0.0000 463.0800 0.1170 ;
      RECT 466.6800 0.0000 487.3940 0.1170 ;
      RECT 490.9940 0.0000 511.3940 0.1170 ;
      RECT 514.9940 0.0000 535.3940 0.1170 ;
      RECT 538.9940 0.0000 559.3940 0.1170 ;
      RECT 562.9940 0.0000 583.3940 0.1170 ;
      RECT 586.9940 0.0000 607.3940 0.1170 ;
      RECT 610.9940 0.0000 631.3940 0.1170 ;
      RECT 634.9940 0.0000 655.3940 0.1170 ;
      RECT 658.9940 0.0000 679.7040 0.1170 ;
      RECT 683.3040 0.0000 704.0140 0.1170 ;
      RECT 707.6140 0.0000 728.3240 0.1170 ;
      RECT 731.9240 0.0000 752.6340 0.1170 ;
      RECT 756.2340 0.0000 776.9440 0.1170 ;
      RECT 780.5440 0.0000 801.2540 0.1170 ;
      RECT 804.8540 0.0000 825.5640 0.1170 ;
      RECT 829.1640 0.0000 849.8740 0.1170 ;
      RECT 853.4740 0.0000 874.1840 0.1170 ;
      RECT 877.7840 0.0000 898.4980 0.1170 ;
      RECT 902.0980 0.0000 922.4980 0.1170 ;
      RECT 926.0980 0.0000 946.4980 0.1170 ;
      RECT 950.0980 0.0000 970.4980 0.1170 ;
      RECT 974.0980 0.0000 994.4980 0.1170 ;
      RECT 998.0980 0.0000 1018.4980 0.1170 ;
      RECT 1022.0980 0.0000 1042.4980 0.1170 ;
      RECT 1046.0980 0.0000 1066.4980 0.1170 ;
      RECT 1070.0980 0.0000 1090.8080 0.1170 ;
      RECT 1094.4080 0.0000 1115.1180 0.1170 ;
      RECT 1118.7180 0.0000 1139.4280 0.1170 ;
      RECT 1143.0280 0.0000 1163.7380 0.1170 ;
      RECT 1167.3380 0.0000 1188.0480 0.1170 ;
      RECT 1191.6480 0.0000 1212.3580 0.1170 ;
      RECT 1215.9580 0.0000 1236.6680 0.1170 ;
      RECT 1240.2680 0.0000 1260.9780 0.1170 ;
      RECT 1264.5780 0.0000 1285.2880 0.1170 ;
      RECT 1288.8880 0.0000 1309.6020 0.1170 ;
      RECT 1313.2020 0.0000 1333.6020 0.1170 ;
      RECT 1337.2020 0.0000 1357.6020 0.1170 ;
      RECT 1361.2020 0.0000 1381.6020 0.1170 ;
      RECT 1385.2020 0.0000 1405.6020 0.1170 ;
      RECT 1409.2020 0.0000 1429.6020 0.1170 ;
      RECT 1433.2020 0.0000 1453.6020 0.1170 ;
      RECT 1457.2020 0.0000 1477.6020 0.1170 ;
      RECT 1481.2020 0.0000 1501.9120 0.1170 ;
      RECT 1505.5120 0.0000 1526.2220 0.1170 ;
      RECT 1529.8220 0.0000 1550.5320 0.1170 ;
      RECT 1554.1320 0.0000 1574.8420 0.1170 ;
      RECT 1578.4420 0.0000 1599.1520 0.1170 ;
      RECT 1602.7520 0.0000 1623.4620 0.1170 ;
      RECT 1627.0620 0.0000 1647.7720 0.1170 ;
      RECT 1651.3720 0.0000 1672.0820 0.1170 ;
      RECT 1675.6820 0.0000 1696.3920 0.1170 ;
      RECT 1699.9920 0.0000 1704.3000 0.1170 ;
      RECT 0.0000 0.1170 1704.3000 640.6830 ;
      RECT 6.9560 640.6830 27.6660 640.8000 ;
      RECT 0.0000 640.6830 3.3560 640.8000 ;
      RECT 31.2660 640.6830 51.9760 640.8000 ;
      RECT 55.5760 640.6830 76.2900 640.8000 ;
      RECT 79.8900 640.6830 100.2900 640.8000 ;
      RECT 103.8900 640.6830 124.2900 640.8000 ;
      RECT 127.8900 640.6830 148.2900 640.8000 ;
      RECT 151.8900 640.6830 172.2900 640.8000 ;
      RECT 175.8900 640.6830 196.2900 640.8000 ;
      RECT 199.8900 640.6830 220.2900 640.8000 ;
      RECT 223.8900 640.6830 244.2900 640.8000 ;
      RECT 247.8900 640.6830 268.6000 640.8000 ;
      RECT 272.2000 640.6830 292.9100 640.8000 ;
      RECT 296.5100 640.6830 317.2200 640.8000 ;
      RECT 320.8200 640.6830 341.5300 640.8000 ;
      RECT 345.1300 640.6830 365.8400 640.8000 ;
      RECT 369.4400 640.6830 390.1500 640.8000 ;
      RECT 393.7500 640.6830 414.4600 640.8000 ;
      RECT 418.0600 640.6830 438.7700 640.8000 ;
      RECT 442.3700 640.6830 463.0800 640.8000 ;
      RECT 466.6800 640.6830 487.3940 640.8000 ;
      RECT 490.9940 640.6830 511.3940 640.8000 ;
      RECT 514.9940 640.6830 535.3940 640.8000 ;
      RECT 538.9940 640.6830 559.3940 640.8000 ;
      RECT 562.9940 640.6830 583.3940 640.8000 ;
      RECT 586.9940 640.6830 607.3940 640.8000 ;
      RECT 610.9940 640.6830 631.3940 640.8000 ;
      RECT 634.9940 640.6830 655.3940 640.8000 ;
      RECT 658.9940 640.6830 679.7040 640.8000 ;
      RECT 683.3040 640.6830 704.0140 640.8000 ;
      RECT 707.6140 640.6830 728.3240 640.8000 ;
      RECT 731.9240 640.6830 752.6340 640.8000 ;
      RECT 756.2340 640.6830 776.9440 640.8000 ;
      RECT 780.5440 640.6830 801.2540 640.8000 ;
      RECT 804.8540 640.6830 825.5640 640.8000 ;
      RECT 829.1640 640.6830 849.8740 640.8000 ;
      RECT 853.4740 640.6830 874.1840 640.8000 ;
      RECT 877.7840 640.6830 898.4980 640.8000 ;
      RECT 902.0980 640.6830 922.4980 640.8000 ;
      RECT 926.0980 640.6830 946.4980 640.8000 ;
      RECT 950.0980 640.6830 970.4980 640.8000 ;
      RECT 974.0980 640.6830 994.4980 640.8000 ;
      RECT 998.0980 640.6830 1018.4980 640.8000 ;
      RECT 1022.0980 640.6830 1042.4980 640.8000 ;
      RECT 1046.0980 640.6830 1066.4980 640.8000 ;
      RECT 1070.0980 640.6830 1090.8080 640.8000 ;
      RECT 1094.4080 640.6830 1115.1180 640.8000 ;
      RECT 1118.7180 640.6830 1139.4280 640.8000 ;
      RECT 1143.0280 640.6830 1163.7380 640.8000 ;
      RECT 1167.3380 640.6830 1188.0480 640.8000 ;
      RECT 1191.6480 640.6830 1212.3580 640.8000 ;
      RECT 1215.9580 640.6830 1236.6680 640.8000 ;
      RECT 1240.2680 640.6830 1260.9780 640.8000 ;
      RECT 1264.5780 640.6830 1285.2880 640.8000 ;
      RECT 1288.8880 640.6830 1309.6020 640.8000 ;
      RECT 1313.2020 640.6830 1333.6020 640.8000 ;
      RECT 1337.2020 640.6830 1357.6020 640.8000 ;
      RECT 1361.2020 640.6830 1381.6020 640.8000 ;
      RECT 1385.2020 640.6830 1405.6020 640.8000 ;
      RECT 1409.2020 640.6830 1429.6020 640.8000 ;
      RECT 1433.2020 640.6830 1453.6020 640.8000 ;
      RECT 1457.2020 640.6830 1477.6020 640.8000 ;
      RECT 1481.2020 640.6830 1501.9120 640.8000 ;
      RECT 1505.5120 640.6830 1526.2220 640.8000 ;
      RECT 1529.8220 640.6830 1550.5320 640.8000 ;
      RECT 1554.1320 640.6830 1574.8420 640.8000 ;
      RECT 1578.4420 640.6830 1599.1520 640.8000 ;
      RECT 1602.7520 640.6830 1623.4620 640.8000 ;
      RECT 1627.0620 640.6830 1647.7720 640.8000 ;
      RECT 1651.3720 640.6830 1672.0820 640.8000 ;
      RECT 1675.6820 640.6830 1696.3920 640.8000 ;
      RECT 1699.9920 640.6830 1704.3000 640.8000 ;
    LAYER M3 ;
      RECT 6.9560 0.0000 27.6660 0.1170 ;
      RECT 0.0000 0.0000 3.3560 0.1170 ;
      RECT 31.2660 0.0000 51.9760 0.1170 ;
      RECT 55.5760 0.0000 76.2900 0.1170 ;
      RECT 79.8900 0.0000 100.2900 0.1170 ;
      RECT 103.8900 0.0000 124.2900 0.1170 ;
      RECT 127.8900 0.0000 148.2900 0.1170 ;
      RECT 151.8900 0.0000 172.2900 0.1170 ;
      RECT 175.8900 0.0000 196.2900 0.1170 ;
      RECT 199.8900 0.0000 220.2900 0.1170 ;
      RECT 223.8900 0.0000 244.2900 0.1170 ;
      RECT 247.8900 0.0000 268.6000 0.1170 ;
      RECT 272.2000 0.0000 292.9100 0.1170 ;
      RECT 296.5100 0.0000 317.2200 0.1170 ;
      RECT 320.8200 0.0000 341.5300 0.1170 ;
      RECT 345.1300 0.0000 365.8400 0.1170 ;
      RECT 369.4400 0.0000 390.1500 0.1170 ;
      RECT 393.7500 0.0000 414.4600 0.1170 ;
      RECT 418.0600 0.0000 438.7700 0.1170 ;
      RECT 442.3700 0.0000 463.0800 0.1170 ;
      RECT 466.6800 0.0000 487.3940 0.1170 ;
      RECT 490.9940 0.0000 511.3940 0.1170 ;
      RECT 514.9940 0.0000 535.3940 0.1170 ;
      RECT 538.9940 0.0000 559.3940 0.1170 ;
      RECT 562.9940 0.0000 583.3940 0.1170 ;
      RECT 586.9940 0.0000 607.3940 0.1170 ;
      RECT 610.9940 0.0000 631.3940 0.1170 ;
      RECT 634.9940 0.0000 655.3940 0.1170 ;
      RECT 658.9940 0.0000 679.7040 0.1170 ;
      RECT 683.3040 0.0000 704.0140 0.1170 ;
      RECT 707.6140 0.0000 728.3240 0.1170 ;
      RECT 731.9240 0.0000 752.6340 0.1170 ;
      RECT 756.2340 0.0000 776.9440 0.1170 ;
      RECT 780.5440 0.0000 801.2540 0.1170 ;
      RECT 804.8540 0.0000 825.5640 0.1170 ;
      RECT 829.1640 0.0000 849.8740 0.1170 ;
      RECT 853.4740 0.0000 874.1840 0.1170 ;
      RECT 877.7840 0.0000 898.4980 0.1170 ;
      RECT 902.0980 0.0000 922.4980 0.1170 ;
      RECT 926.0980 0.0000 946.4980 0.1170 ;
      RECT 950.0980 0.0000 970.4980 0.1170 ;
      RECT 974.0980 0.0000 994.4980 0.1170 ;
      RECT 998.0980 0.0000 1018.4980 0.1170 ;
      RECT 1022.0980 0.0000 1042.4980 0.1170 ;
      RECT 1046.0980 0.0000 1066.4980 0.1170 ;
      RECT 1070.0980 0.0000 1090.8080 0.1170 ;
      RECT 1094.4080 0.0000 1115.1180 0.1170 ;
      RECT 1118.7180 0.0000 1139.4280 0.1170 ;
      RECT 1143.0280 0.0000 1163.7380 0.1170 ;
      RECT 1167.3380 0.0000 1188.0480 0.1170 ;
      RECT 1191.6480 0.0000 1212.3580 0.1170 ;
      RECT 1215.9580 0.0000 1236.6680 0.1170 ;
      RECT 1240.2680 0.0000 1260.9780 0.1170 ;
      RECT 1264.5780 0.0000 1285.2880 0.1170 ;
      RECT 1288.8880 0.0000 1309.6020 0.1170 ;
      RECT 1313.2020 0.0000 1333.6020 0.1170 ;
      RECT 1337.2020 0.0000 1357.6020 0.1170 ;
      RECT 1361.2020 0.0000 1381.6020 0.1170 ;
      RECT 1385.2020 0.0000 1405.6020 0.1170 ;
      RECT 1409.2020 0.0000 1429.6020 0.1170 ;
      RECT 1433.2020 0.0000 1453.6020 0.1170 ;
      RECT 1457.2020 0.0000 1477.6020 0.1170 ;
      RECT 1481.2020 0.0000 1501.9120 0.1170 ;
      RECT 1505.5120 0.0000 1526.2220 0.1170 ;
      RECT 1529.8220 0.0000 1550.5320 0.1170 ;
      RECT 1554.1320 0.0000 1574.8420 0.1170 ;
      RECT 1578.4420 0.0000 1599.1520 0.1170 ;
      RECT 1602.7520 0.0000 1623.4620 0.1170 ;
      RECT 1627.0620 0.0000 1647.7720 0.1170 ;
      RECT 1651.3720 0.0000 1672.0820 0.1170 ;
      RECT 1675.6820 0.0000 1696.3920 0.1170 ;
      RECT 1699.9920 0.0000 1704.3000 0.1170 ;
      RECT 0.0000 0.1170 1704.3000 640.6830 ;
      RECT 6.9560 640.6830 27.6660 640.8000 ;
      RECT 0.0000 640.6830 3.3560 640.8000 ;
      RECT 31.2660 640.6830 51.9760 640.8000 ;
      RECT 55.5760 640.6830 76.2900 640.8000 ;
      RECT 79.8900 640.6830 100.2900 640.8000 ;
      RECT 103.8900 640.6830 124.2900 640.8000 ;
      RECT 127.8900 640.6830 148.2900 640.8000 ;
      RECT 151.8900 640.6830 172.2900 640.8000 ;
      RECT 175.8900 640.6830 196.2900 640.8000 ;
      RECT 199.8900 640.6830 220.2900 640.8000 ;
      RECT 223.8900 640.6830 244.2900 640.8000 ;
      RECT 247.8900 640.6830 268.6000 640.8000 ;
      RECT 272.2000 640.6830 292.9100 640.8000 ;
      RECT 296.5100 640.6830 317.2200 640.8000 ;
      RECT 320.8200 640.6830 341.5300 640.8000 ;
      RECT 345.1300 640.6830 365.8400 640.8000 ;
      RECT 369.4400 640.6830 390.1500 640.8000 ;
      RECT 393.7500 640.6830 414.4600 640.8000 ;
      RECT 418.0600 640.6830 438.7700 640.8000 ;
      RECT 442.3700 640.6830 463.0800 640.8000 ;
      RECT 466.6800 640.6830 487.3940 640.8000 ;
      RECT 490.9940 640.6830 511.3940 640.8000 ;
      RECT 514.9940 640.6830 535.3940 640.8000 ;
      RECT 538.9940 640.6830 559.3940 640.8000 ;
      RECT 562.9940 640.6830 583.3940 640.8000 ;
      RECT 586.9940 640.6830 607.3940 640.8000 ;
      RECT 610.9940 640.6830 631.3940 640.8000 ;
      RECT 634.9940 640.6830 655.3940 640.8000 ;
      RECT 658.9940 640.6830 679.7040 640.8000 ;
      RECT 683.3040 640.6830 704.0140 640.8000 ;
      RECT 707.6140 640.6830 728.3240 640.8000 ;
      RECT 731.9240 640.6830 752.6340 640.8000 ;
      RECT 756.2340 640.6830 776.9440 640.8000 ;
      RECT 780.5440 640.6830 801.2540 640.8000 ;
      RECT 804.8540 640.6830 825.5640 640.8000 ;
      RECT 829.1640 640.6830 849.8740 640.8000 ;
      RECT 853.4740 640.6830 874.1840 640.8000 ;
      RECT 877.7840 640.6830 898.4980 640.8000 ;
      RECT 902.0980 640.6830 922.4980 640.8000 ;
      RECT 926.0980 640.6830 946.4980 640.8000 ;
      RECT 950.0980 640.6830 970.4980 640.8000 ;
      RECT 974.0980 640.6830 994.4980 640.8000 ;
      RECT 998.0980 640.6830 1018.4980 640.8000 ;
      RECT 1022.0980 640.6830 1042.4980 640.8000 ;
      RECT 1046.0980 640.6830 1066.4980 640.8000 ;
      RECT 1070.0980 640.6830 1090.8080 640.8000 ;
      RECT 1094.4080 640.6830 1115.1180 640.8000 ;
      RECT 1118.7180 640.6830 1139.4280 640.8000 ;
      RECT 1143.0280 640.6830 1163.7380 640.8000 ;
      RECT 1167.3380 640.6830 1188.0480 640.8000 ;
      RECT 1191.6480 640.6830 1212.3580 640.8000 ;
      RECT 1215.9580 640.6830 1236.6680 640.8000 ;
      RECT 1240.2680 640.6830 1260.9780 640.8000 ;
      RECT 1264.5780 640.6830 1285.2880 640.8000 ;
      RECT 1288.8880 640.6830 1309.6020 640.8000 ;
      RECT 1313.2020 640.6830 1333.6020 640.8000 ;
      RECT 1337.2020 640.6830 1357.6020 640.8000 ;
      RECT 1361.2020 640.6830 1381.6020 640.8000 ;
      RECT 1385.2020 640.6830 1405.6020 640.8000 ;
      RECT 1409.2020 640.6830 1429.6020 640.8000 ;
      RECT 1433.2020 640.6830 1453.6020 640.8000 ;
      RECT 1457.2020 640.6830 1477.6020 640.8000 ;
      RECT 1481.2020 640.6830 1501.9120 640.8000 ;
      RECT 1505.5120 640.6830 1526.2220 640.8000 ;
      RECT 1529.8220 640.6830 1550.5320 640.8000 ;
      RECT 1554.1320 640.6830 1574.8420 640.8000 ;
      RECT 1578.4420 640.6830 1599.1520 640.8000 ;
      RECT 1602.7520 640.6830 1623.4620 640.8000 ;
      RECT 1627.0620 640.6830 1647.7720 640.8000 ;
      RECT 1651.3720 640.6830 1672.0820 640.8000 ;
      RECT 1675.6820 640.6830 1696.3920 640.8000 ;
      RECT 1699.9920 640.6830 1704.3000 640.8000 ;
    LAYER M2 ;
      RECT 0.0000 0.2770 1704.3000 640.5230 ;
    LAYER M1 ;
      RECT 0.0000 0.0000 1704.3000 640.8000 ;
  END
END fe

END LIBRARY
