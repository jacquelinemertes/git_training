module fft512_tb #(
	parameter NBW_IN    = 'd9,
    parameter NBI_IN    = 'd2,
    parameter NBW_OUT   = NBW_IN,
    parameter NBI_OUT   = NBI_IN,
	parameter NBW_FFT   = NBW_IN+5,
    parameter NBI_FFT   = NBI_IN+5
)
( );
	logic clk;
    logic rst_async_n;  

    logic i_valid;

  	logic signed [NBW_IN-1:0] i_data_i [0:63];
    logic signed [NBW_IN-1:0] i_data_q [0:63];

	logic o_valid_hi, o_valid_lo;			
	
    logic signed [NBW_FFT-1:0] o_data_lo_i [0:63];
    logic signed [NBW_FFT-1:0] o_data_lo_q [0:63];
	logic signed [NBW_FFT-1:0] o_data_hi_i [0:63];
    logic signed [NBW_FFT-1:0] o_data_hi_q [0:63];

integer j;

fft512 #(
        .NBW_IN (NBW_IN ),
        .NBI_IN (NBI_IN ),
        .NBW_OUT(NBW_FFT),
        .NBI_OUT(NBI_FFT)
    ) uu_fft512
    (   
        .clk        (clk        ),
        .rst_async_n(rst_async_n),
        .i_overlap  (0  ),
        .i_valid    (i_valid    ),
        .i_data_i   (i_data_i   ),
        .i_data_q   (i_data_q   ),

        .o_valid_lo (o_valid_lo ),
        .o_data_lo_i(o_data_lo_i),
        .o_data_lo_q(o_data_lo_q),

        .o_valid_hi (o_valid_hi ),
        .o_data_hi_i(o_data_hi_i),
        .o_data_hi_q(o_data_hi_q)
    );
always begin
	#1
	clk = ~clk;
end

initial begin
	clk = 0;
	rst_async_n = 0;
	i_valid = 0;
	#5
	rst_async_n = 1;
	#2
i_valid = 1;
/*i_data_i[0] = 9'd114;		//sample 0
i_data_q[0] =-9'd43;
i_data_i[1] = 9'd90;		//sample 1
i_data_q[1] = 9'd41;
i_data_i[2] = 9'd50;		//sample 2
i_data_q[2] =-9'd94;
i_data_i[3] =-9'd112;		//sample 3
i_data_q[3] = 9'd52;
i_data_i[4] = 9'd26;		//sample 4
i_data_q[4] =-9'd14;
i_data_i[5] =-9'd76;		//sample 5
i_data_q[5] =-9'd38;
i_data_i[6] =-9'd8;			//sample 6
i_data_q[6] =-9'd150;
i_data_i[7] = 9'd17;		//sample 7
i_data_q[7] =-9'd125;
i_data_i[8] = 9'd114;		//sample 8
i_data_q[8] = 9'd29;
i_data_i[9] = 9'd56;		//sample 9
i_data_q[9] = 9'd85;
i_data_i[10] =-9'd76;		//sample 10
i_data_q[10] = 9'd7;
i_data_i[11] =-9'd42;		//sample 11
i_data_q[11] = 9'd44;
i_data_i[12] = 9'd36;		//sample 12
i_data_q[12] = 9'd110;
i_data_i[13] = 9'd16;		//sample 13
i_data_q[13] = 9'd90;
i_data_i[14] =-9'd28;		//sample 14
i_data_q[14] = 9'd76;
i_data_i[15] =-9'd4;		//sample 15
i_data_q[15] =-9'd98;
i_data_i[16] = 9'd125;		//sample 16
i_data_q[16] =-9'd38;
i_data_i[17] =-9'd33;		//sample 17
i_data_q[17] = 9'd11;
i_data_i[18] =-9'd84;		//sample 18
i_data_q[18] = 9'd50;
i_data_i[19] =-9'd67;		//sample 19
i_data_q[19] =-9'd94;
i_data_i[20] =-9'd36;		//sample 20
i_data_q[20] =-9'd0;
i_data_i[21] = 9'd73;		//sample 21
i_data_q[21] = 9'd58;
i_data_i[22] =-9'd118;		//sample 22
i_data_q[22] =-9'd49;
i_data_i[23] =-9'd106;		//sample 23
i_data_q[23] =-9'd89;
i_data_i[24] = 9'd33;		//sample 24
i_data_q[24] = 9'd114;
i_data_i[25] =-9'd32;		//sample 25
i_data_q[25] = 9'd21;
i_data_i[26] = 9'd90;		//sample 26
i_data_q[26] =-9'd32;
i_data_i[27] = 9'd62;		//sample 27
i_data_q[27] = 9'd123;
i_data_i[28] =-9'd114;		//sample 28
i_data_q[28] = 9'd68;
i_data_i[29] =-9'd34;		//sample 29
i_data_q[29] =-9'd121;
i_data_i[30] = 9'd16;		//sample 30
i_data_q[30] = 9'd146;
i_data_i[31] =-9'd98;		//sample 31
i_data_q[31] = 9'd47;
i_data_i[32] = 9'd49;		//sample 32
i_data_q[32] = 9'd22;
i_data_i[33] =-9'd102;		//sample 33
i_data_q[33] = 9'd5;
i_data_i[34] =-9'd115;		//sample 34
i_data_q[34] =-9'd57;
i_data_i[35] =-9'd45;		//sample 35
i_data_q[35] = 9'd3;
i_data_i[36] =-9'd26;		//sample 36
i_data_q[36] = 9'd48;
i_data_i[37] =-9'd76;		//sample 37
i_data_q[37] = 9'd49;
i_data_i[38] =-9'd104;		//sample 38
i_data_q[38] =-9'd122;
i_data_i[39] = 9'd25;		//sample 39
i_data_q[39] =-9'd28;
i_data_i[40] =-9'd67;		//sample 40
i_data_q[40] = 9'd90;
i_data_i[41] = 9'd54;		//sample 41
i_data_q[41] =-9'd87;
i_data_i[42] = 9'd58;		//sample 42
i_data_q[42] = 9'd83;
i_data_i[43] = 9'd6;		//sample 43
i_data_q[43] =-9'd52;
i_data_i[44] =-9'd1;		//sample 44
i_data_q[44] = 9'd37;
i_data_i[45] =-9'd44;		//sample 45
i_data_q[45] = 9'd69;
i_data_i[46] =-9'd87;		//sample 46
i_data_q[46] = 9'd70;
i_data_i[47] =-9'd32;		//sample 47
i_data_q[47] =-9'd7;
i_data_i[48] = 9'd74;		//sample 48
i_data_q[48] =-9'd112;
i_data_i[49] = 9'd43;		//sample 49
i_data_q[49] =-9'd39;
i_data_i[50] =-9'd105;		//sample 50
i_data_q[50] = 9'd84;
i_data_i[51] =-9'd82;		//sample 51
i_data_q[51] =-9'd112;
i_data_i[52] =-9'd87;		//sample 52
i_data_q[52] =-9'd35;
i_data_i[53] =-9'd5;		//sample 53
i_data_q[53] =-9'd54;
i_data_i[54] =-9'd26;		//sample 54
i_data_q[54] =-9'd45;
i_data_i[55] = 9'd81;		//sample 55
i_data_q[55] =-9'd37;
i_data_i[56] = 9'd55;		//sample 56
i_data_q[56] =-9'd9;
i_data_i[57] = 9'd65;		//sample 57
i_data_q[57] = 9'd98;
i_data_i[58] =-9'd70;		//sample 58
i_data_q[58] =-9'd88;
i_data_i[59] = 9'd83;		//sample 59
i_data_q[59] = 9'd53;
i_data_i[60] =-9'd93;		//sample 60
i_data_q[60] =-9'd2;
i_data_i[61] =-9'd24;		//sample 61
i_data_q[61] = 9'd45;
i_data_i[62] = 9'd25;		//sample 62
i_data_q[62] =-9'd26;
i_data_i[63] = 9'd27;		//sample 63
i_data_q[63] = 9'd101;
#2
i_data_i[0] = 9'd8;		//sample 64
i_data_q[0] = 9'd82;
i_data_i[1] =-9'd6;		//sample 65
i_data_q[1] =-9'd30;
i_data_i[2] = 9'd102;		//sample 66
i_data_q[2] =-9'd36;
i_data_i[3] = 9'd30;		//sample 67
i_data_q[3] = 9'd36;
i_data_i[4] = 9'd92;		//sample 68
i_data_q[4] = 9'd18;
i_data_i[5] = 9'd6;		//sample 69
i_data_q[5] =-9'd162;
i_data_i[6] =-9'd17;		//sample 70
i_data_q[6] = 9'd116;
i_data_i[7] =-9'd106;		//sample 71
i_data_q[7] = 9'd14;
i_data_i[8] =-9'd42;		//sample 72
i_data_q[8] = 9'd118;
i_data_i[9] = 9'd121;		//sample 73
i_data_q[9] = 9'd67;
i_data_i[10] = 9'd111;		//sample 74
i_data_q[10] = 9'd8;
i_data_i[11] =-9'd93;		//sample 75
i_data_q[11] =-9'd18;
i_data_i[12] = 9'd101;		//sample 76
i_data_q[12] = 9'd124;
i_data_i[13] = 9'd9;		//sample 77
i_data_q[13] = 9'd116;
i_data_i[14] = 9'd35;		//sample 78
i_data_q[14] =-9'd10;
i_data_i[15] = 9'd28;		//sample 79
i_data_q[15] =-9'd19;
i_data_i[16] =-9'd56;		//sample 80
i_data_q[16] =-9'd61;
i_data_i[17] =-9'd19;		//sample 81
i_data_q[17] = 9'd142;
i_data_i[18] = 9'd73;		//sample 82
i_data_q[18] = 9'd68;
i_data_i[19] =-9'd89;		//sample 83
i_data_q[19] =-9'd49;
i_data_i[20] =-9'd129;		//sample 84
i_data_q[20] =-9'd57;
i_data_i[21] = 9'd130;		//sample 85
i_data_q[21] = 9'd81;
i_data_i[22] =-9'd89;		//sample 86
i_data_q[22] =-9'd13;
i_data_i[23] = 9'd47;		//sample 87
i_data_q[23] = 9'd84;
i_data_i[24] = 9'd90;		//sample 88
i_data_q[24] =-9'd95;
i_data_i[25] = 9'd97;		//sample 89
i_data_q[25] = 9'd63;
i_data_i[26] =-9'd105;		//sample 90
i_data_q[26] = 9'd47;
i_data_i[27] = 9'd69;		//sample 91
i_data_q[27] =-9'd23;
i_data_i[28] = 9'd151;		//sample 92
i_data_q[28] =-9'd38;
i_data_i[29] = 9'd69;		//sample 93
i_data_q[29] = 9'd76;
i_data_i[30] =-9'd90;		//sample 94
i_data_q[30] = 9'd58;
i_data_i[31] =-9'd40;		//sample 95
i_data_q[31] =-9'd100;
i_data_i[32] =-9'd105;		//sample 96
i_data_q[32] =-9'd34;
i_data_i[33] = 9'd54;		//sample 97
i_data_q[33] =-9'd119;
i_data_i[34] =-9'd19;		//sample 98
i_data_q[34] = 9'd18;
i_data_i[35] =-9'd106;		//sample 99
i_data_q[35] =-9'd8;
i_data_i[36] =-9'd29;		//sample 100
i_data_q[36] =-9'd79;
i_data_i[37] =-9'd104;		//sample 101
i_data_q[37] = 9'd69;
i_data_i[38] =-9'd1;		//sample 102
i_data_q[38] = 9'd53;
i_data_i[39] = 9'd37;		//sample 103
i_data_q[39] =-9'd1;
i_data_i[40] =-9'd42;		//sample 104
i_data_q[40] = 9'd101;
i_data_i[41] = 9'd2;		//sample 105
i_data_q[41] =-9'd59;
i_data_i[42] = 9'd35;		//sample 106
i_data_q[42] = 9'd0;
i_data_i[43] = 9'd58;		//sample 107
i_data_q[43] =-9'd64;
i_data_i[44] = 9'd70;		//sample 108
i_data_q[44] = 9'd88;
i_data_i[45] =-9'd76;		//sample 109
i_data_q[45] = 9'd64;
i_data_i[46] =-9'd101;		//sample 110
i_data_q[46] = 9'd57;
i_data_i[47] =-9'd97;		//sample 111
i_data_q[47] = 9'd2;
i_data_i[48] =-9'd99;		//sample 112
i_data_q[48] =-9'd87;
i_data_i[49] = 9'd16;		//sample 113
i_data_q[49] = 9'd40;
i_data_i[50] =-9'd76;		//sample 114
i_data_q[50] =-9'd64;
i_data_i[51] =-9'd35;		//sample 115
i_data_q[51] = 9'd25;
i_data_i[52] = 9'd36;		//sample 116
i_data_q[52] = 9'd119;
i_data_i[53] = 9'd44;		//sample 117
i_data_q[53] = 9'd6;
i_data_i[54] =-9'd82;		//sample 118
i_data_q[54] =-9'd32;
i_data_i[55] = 9'd111;		//sample 119
i_data_q[55] =-9'd46;
i_data_i[56] =-9'd0;		//sample 120
i_data_q[56] =-9'd57;
i_data_i[57] = 9'd31;		//sample 121
i_data_q[57] = 9'd81;
i_data_i[58] = 9'd89;		//sample 122
i_data_q[58] =-9'd76;
i_data_i[59] = 9'd30;		//sample 123
i_data_q[59] = 9'd14;
i_data_i[60] =-9'd19;		//sample 124
i_data_q[60] = 9'd108;
i_data_i[61] = 9'd88;		//sample 125
i_data_q[61] = 9'd83;
i_data_i[62] = 9'd109;		//sample 126
i_data_q[62] =-9'd34;
i_data_i[63] =-9'd2;		//sample 127
i_data_q[63] =-9'd100;
#2
i_data_i[0] = 9'd48;		//sample 128
i_data_q[0] =-9'd10;
i_data_i[1] =-9'd76;		//sample 129
i_data_q[1] =-9'd95;
i_data_i[2] =-9'd9;		//sample 130
i_data_q[2] =-9'd136;
i_data_i[3] =-9'd43;		//sample 131
i_data_q[3] =-9'd16;
i_data_i[4] = 9'd16;		//sample 132
i_data_q[4] = 9'd98;
i_data_i[5] =-9'd31;		//sample 133
i_data_q[5] = 9'd124;
i_data_i[6] = 9'd62;		//sample 134
i_data_q[6] =-9'd112;
i_data_i[7] = 9'd15;		//sample 135
i_data_q[7] =-9'd104;
i_data_i[8] = 9'd11;		//sample 136
i_data_q[8] =-9'd89;
i_data_i[9] =-9'd83;		//sample 137
i_data_q[9] =-9'd18;
i_data_i[10] =-9'd115;		//sample 138
i_data_q[10] = 9'd85;
i_data_i[11] =-9'd76;		//sample 139
i_data_q[11] =-9'd94;
i_data_i[12] = 9'd1;		//sample 140
i_data_q[12] =-9'd46;
i_data_i[13] = 9'd116;		//sample 141
i_data_q[13] =-9'd71;
i_data_i[14] =-9'd73;		//sample 142
i_data_q[14] = 9'd65;
i_data_i[15] =-9'd102;		//sample 143
i_data_q[15] = 9'd40;
i_data_i[16] =-9'd24;		//sample 144
i_data_q[16] = 9'd7;
i_data_i[17] = 9'd45;		//sample 145
i_data_q[17] = 9'd5;
i_data_i[18] =-9'd63;		//sample 146
i_data_q[18] =-9'd13;
i_data_i[19] =-9'd1;		//sample 147
i_data_q[19] =-9'd42;
i_data_i[20] =-9'd31;		//sample 148
i_data_q[20] =-9'd37;
i_data_i[21] = 9'd9;		//sample 149
i_data_q[21] =-9'd92;
i_data_i[22] =-9'd35;		//sample 150
i_data_q[22] =-9'd26;
i_data_i[23] =-9'd91;		//sample 151
i_data_q[23] =-9'd111;
i_data_i[24] = 9'd125;		//sample 152
i_data_q[24] =-9'd66;
i_data_i[25] = 9'd13;		//sample 153
i_data_q[25] = 9'd98;
i_data_i[26] =-9'd27;		//sample 154
i_data_q[26] = 9'd25;
i_data_i[27] = 9'd42;		//sample 155
i_data_q[27] =-9'd93;
i_data_i[28] =-9'd56;		//sample 156
i_data_q[28] =-9'd2;
i_data_i[29] = 9'd71;		//sample 157
i_data_q[29] = 9'd44;
i_data_i[30] = 9'd26;		//sample 158
i_data_q[30] =-9'd130;
i_data_i[31] =-9'd47;		//sample 159
i_data_q[31] = 9'd152;
i_data_i[32] = 9'd112;		//sample 160
i_data_q[32] = 9'd17;
i_data_i[33] = 9'd9;		//sample 161
i_data_q[33] =-9'd55;
i_data_i[34] = 9'd22;		//sample 162
i_data_q[34] =-9'd108;
i_data_i[35] =-9'd28;		//sample 163
i_data_q[35] = 9'd111;
i_data_i[36] =-9'd3;		//sample 164
i_data_q[36] = 9'd88;
i_data_i[37] = 9'd80;		//sample 165
i_data_q[37] = 9'd4;
i_data_i[38] = 9'd3;		//sample 166
i_data_q[38] =-9'd101;
i_data_i[39] = 9'd57;		//sample 167
i_data_q[39] = 9'd73;
i_data_i[40] =-9'd28;		//sample 168
i_data_q[40] = 9'd16;
i_data_i[41] =-9'd8;		//sample 169
i_data_q[41] =-9'd130;
i_data_i[42] = 9'd33;		//sample 170
i_data_q[42] =-9'd119;
i_data_i[43] = 9'd87;		//sample 171
i_data_q[43] = 9'd65;
i_data_i[44] = 9'd7;		//sample 172
i_data_q[44] = 9'd105;
i_data_i[45] =-9'd97;		//sample 173
i_data_q[45] = 9'd38;
i_data_i[46] =-9'd29;		//sample 174
i_data_q[46] = 9'd57;
i_data_i[47] =-9'd39;		//sample 175
i_data_q[47] =-9'd80;
i_data_i[48] = 9'd81;		//sample 176
i_data_q[48] = 9'd111;
i_data_i[49] =-9'd59;		//sample 177
i_data_q[49] = 9'd83;
i_data_i[50] = 9'd83;		//sample 178
i_data_q[50] =-9'd2;
i_data_i[51] =-9'd31;		//sample 179
i_data_q[51] = 9'd109;
i_data_i[52] = 9'd73;		//sample 180
i_data_q[52] = 9'd76;
i_data_i[53] = 9'd35;		//sample 181
i_data_q[53] =-9'd18;
i_data_i[54] = 9'd32;		//sample 182
i_data_q[54] = 9'd100;
i_data_i[55] =-9'd136;		//sample 183
i_data_q[55] =-9'd43;
i_data_i[56] = 9'd3;		//sample 184
i_data_q[56] = 9'd91;
i_data_i[57] = 9'd22;		//sample 185
i_data_q[57] =-9'd43;
i_data_i[58] = 9'd87;		//sample 186
i_data_q[58] =-9'd52;
i_data_i[59] =-9'd90;		//sample 187
i_data_q[59] = 9'd90;
i_data_i[60] =-9'd31;		//sample 188
i_data_q[60] =-9'd92;
i_data_i[61] = 9'd24;		//sample 189
i_data_q[61] = 9'd48;
i_data_i[62] = 9'd126;		//sample 190
i_data_q[62] =-9'd44;
i_data_i[63] = 9'd87;		//sample 191
i_data_q[63] = 9'd62;
#2
i_data_i[0] = 9'd101;		//sample 192
i_data_q[0] = 9'd41;
i_data_i[1] =-9'd13;		//sample 193
i_data_q[1] =-9'd124;
i_data_i[2] =-9'd8;		//sample 194
i_data_q[2] =-9'd147;
i_data_i[3] =-9'd56;		//sample 195
i_data_q[3] = 9'd12;
i_data_i[4] = 9'd11;		//sample 196
i_data_q[4] = 9'd111;
i_data_i[5] =-9'd34;		//sample 197
i_data_q[5] = 9'd117;
i_data_i[6] = 9'd84;		//sample 198
i_data_q[6] =-9'd141;
i_data_i[7] =-9'd101;		//sample 199
i_data_q[7] = 9'd108;
i_data_i[8] = 9'd33;		//sample 200
i_data_q[8] = 9'd21;
i_data_i[9] =-9'd38;		//sample 201
i_data_q[9] =-9'd43;
i_data_i[10] = 9'd89;		//sample 202
i_data_q[10] =-9'd5;
i_data_i[11] = 9'd83;		//sample 203
i_data_q[11] =-9'd88;
i_data_i[12] =-9'd21;		//sample 204
i_data_q[12] = 9'd106;
i_data_i[13] =-9'd73;		//sample 205
i_data_q[13] =-9'd66;
i_data_i[14] =-9'd96;		//sample 206
i_data_q[14] = 9'd46;
i_data_i[15] =-9'd58;		//sample 207
i_data_q[15] = 9'd4;
i_data_i[16] = 9'd73;		//sample 208
i_data_q[16] = 9'd76;
i_data_i[17] = 9'd71;		//sample 209
i_data_q[17] = 9'd95;
i_data_i[18] =-9'd107;		//sample 210
i_data_q[18] = 9'd15;
i_data_i[19] = 9'd30;		//sample 211
i_data_q[19] =-9'd109;
i_data_i[20] =-9'd119;		//sample 212
i_data_q[20] =-9'd105;
i_data_i[21] = 9'd56;		//sample 213
i_data_q[21] =-9'd100;
i_data_i[22] = 9'd4;		//sample 214
i_data_q[22] = 9'd34;
i_data_i[23] =-9'd81;		//sample 215
i_data_q[23] = 9'd5;
i_data_i[24] = 9'd115;		//sample 216
i_data_q[24] = 9'd3;
i_data_i[25] = 9'd91;		//sample 217
i_data_q[25] =-9'd60;
i_data_i[26] = 9'd1;		//sample 218
i_data_q[26] = 9'd39;
i_data_i[27] = 9'd23;		//sample 219
i_data_q[27] = 9'd92;
i_data_i[28] = 9'd98;		//sample 220
i_data_q[28] =-9'd6;
i_data_i[29] = 9'd91;		//sample 221
i_data_q[29] =-9'd5;
i_data_i[30] = 9'd37;		//sample 222
i_data_q[30] = 9'd38;
i_data_i[31] = 9'd119;		//sample 223
i_data_q[31] = 9'd86;
i_data_i[32] =-9'd14;		//sample 224
i_data_q[32] = 9'd116;
i_data_i[33] = 9'd104;		//sample 225
i_data_q[33] = 9'd106;
i_data_i[34] =-9'd103;		//sample 226
i_data_q[34] = 9'd23;
i_data_i[35] =-9'd110;		//sample 227
i_data_q[35] = 9'd9;
i_data_i[36] = 9'd36;		//sample 228
i_data_q[36] =-9'd10;
i_data_i[37] = 9'd47;		//sample 229
i_data_q[37] = 9'd128;
i_data_i[38] =-9'd50;		//sample 230
i_data_q[38] =-9'd11;
i_data_i[39] =-9'd40;		//sample 231
i_data_q[39] =-9'd75;
i_data_i[40] =-9'd18;		//sample 232
i_data_q[40] = 9'd154;
i_data_i[41] = 9'd63;		//sample 233
i_data_q[41] = 9'd76;
i_data_i[42] =-9'd64;		//sample 234
i_data_q[42] =-9'd19;
i_data_i[43] =-9'd92;		//sample 235
i_data_q[43] = 9'd80;
i_data_i[44] =-9'd44;		//sample 236
i_data_q[44] =-9'd32;
i_data_i[45] = 9'd105;		//sample 237
i_data_q[45] =-9'd22;
i_data_i[46] =-9'd85;		//sample 238
i_data_q[46] =-9'd54;
i_data_i[47] =-9'd74;		//sample 239
i_data_q[47] =-9'd51;
i_data_i[48] =-9'd99;		//sample 240
i_data_q[48] = 9'd8;
i_data_i[49] =-9'd9;		//sample 241
i_data_q[49] =-9'd41;
i_data_i[50] =-9'd100;		//sample 242
i_data_q[50] =-9'd18;
i_data_i[51] = 9'd6;		//sample 243
i_data_q[51] = 9'd119;
i_data_i[52] = 9'd4;		//sample 244
i_data_q[52] =-9'd137;
i_data_i[53] =-9'd24;		//sample 245
i_data_q[53] = 9'd147;
i_data_i[54] =-9'd105;		//sample 246
i_data_q[54] = 9'd8;
i_data_i[55] = 9'd78;		//sample 247
i_data_q[55] =-9'd79;
i_data_i[56] =-9'd95;		//sample 248
i_data_q[56] = 9'd43;
i_data_i[57] = 9'd92;		//sample 249
i_data_q[57] = 9'd7;
i_data_i[58] =-9'd90;		//sample 250
i_data_q[58] = 9'd91;
i_data_i[59] = 9'd119;		//sample 251
i_data_q[59] =-9'd70;
i_data_i[60] =-9'd117;		//sample 252
i_data_q[60] = 9'd50;
i_data_i[61] = 9'd55;		//sample 253
i_data_q[61] = 9'd1;
i_data_i[62] =-9'd65;		//sample 254
i_data_q[62] =-9'd75;
i_data_i[63] =-9'd30;		//sample 255
i_data_q[63] =-9'd156;
#2
i_data_i[0] = 9'd34;		//sample 256
i_data_q[0] = 9'd135;
i_data_i[1] = 9'd13;		//sample 257
i_data_q[1] = 9'd92;
i_data_i[2] =-9'd62;		//sample 258
i_data_q[2] =-9'd58;
i_data_i[3] = 9'd48;		//sample 259
i_data_q[3] = 9'd63;
i_data_i[4] =-9'd21;		//sample 260
i_data_q[4] =-9'd22;
i_data_i[5] = 9'd29;		//sample 261
i_data_q[5] = 9'd6;
i_data_i[6] =-9'd105;		//sample 262
i_data_q[6] = 9'd92;
i_data_i[7] =-9'd18;		//sample 263
i_data_q[7] =-9'd29;
i_data_i[8] =-9'd45;		//sample 264
i_data_q[8] = 9'd38;
i_data_i[9] = 9'd91;		//sample 265
i_data_q[9] = 9'd54;
i_data_i[10] =-9'd48;		//sample 266
i_data_q[10] = 9'd14;
i_data_i[11] =-9'd17;		//sample 267
i_data_q[11] =-9'd59;
i_data_i[12] =-9'd81;		//sample 268
i_data_q[12] =-9'd24;
i_data_i[13] =-9'd43;		//sample 269
i_data_q[13] = 9'd84;
i_data_i[14] = 9'd9;		//sample 270
i_data_q[14] = 9'd87;
i_data_i[15] = 9'd72;		//sample 271
i_data_q[15] = 9'd54;
i_data_i[16] =-9'd83;		//sample 272
i_data_q[16] =-9'd81;
i_data_i[17] =-9'd37;		//sample 273
i_data_q[17] = 9'd44;
i_data_i[18] =-9'd91;		//sample 274
i_data_q[18] = 9'd120;
i_data_i[19] = 9'd107;		//sample 275
i_data_q[19] = 9'd33;
i_data_i[20] = 9'd36;		//sample 276
i_data_q[20] =-9'd73;
i_data_i[21] = 9'd74;		//sample 277
i_data_q[21] = 9'd35;
i_data_i[22] =-9'd142;		//sample 278
i_data_q[22] = 9'd59;
i_data_i[23] = 9'd110;		//sample 279
i_data_q[23] =-9'd29;
i_data_i[24] =-9'd14;		//sample 280
i_data_q[24] = 9'd88;
i_data_i[25] =-9'd94;		//sample 281
i_data_q[25] = 9'd61;
i_data_i[26] = 9'd73;		//sample 282
i_data_q[26] = 9'd41;
i_data_i[27] = 9'd20;		//sample 283
i_data_q[27] =-9'd109;
i_data_i[28] =-9'd56;		//sample 284
i_data_q[28] =-9'd82;
i_data_i[29] = 9'd21;		//sample 285
i_data_q[29] =-9'd18;
i_data_i[30] = 9'd111;		//sample 286
i_data_q[30] = 9'd83;
i_data_i[31] =-9'd52;		//sample 287
i_data_q[31] =-9'd46;
i_data_i[32] =-9'd87;		//sample 288
i_data_q[32] =-9'd93;
i_data_i[33] =-9'd111;		//sample 289
i_data_q[33] = 9'd91;
i_data_i[34] =-9'd114;		//sample 290
i_data_q[34] =-9'd17;
i_data_i[35] =-9'd44;		//sample 291
i_data_q[35] = 9'd3;
i_data_i[36] =-9'd107;		//sample 292
i_data_q[36] = 9'd21;
i_data_i[37] = 9'd86;		//sample 293
i_data_q[37] =-9'd70;
i_data_i[38] = 9'd38;		//sample 294
i_data_q[38] = 9'd117;
i_data_i[39] = 9'd145;		//sample 295
i_data_q[39] = 9'd9;
i_data_i[40] = 9'd84;		//sample 296
i_data_q[40] =-9'd72;
i_data_i[41] = 9'd85;		//sample 297
i_data_q[41] = 9'd3;
i_data_i[42] =-9'd40;		//sample 298
i_data_q[42] = 9'd51;
i_data_i[43] =-9'd66;		//sample 299
i_data_q[43] = 9'd108;
i_data_i[44] =-9'd102;		//sample 300
i_data_q[44] =-9'd48;
i_data_i[45] =-9'd15;		//sample 301
i_data_q[45] =-9'd88;
i_data_i[46] = 9'd107;		//sample 302
i_data_q[46] =-9'd74;
i_data_i[47] =-9'd52;		//sample 303
i_data_q[47] = 9'd79;
i_data_i[48] =-9'd63;		//sample 304
i_data_q[48] = 9'd5;
i_data_i[49] =-9'd134;		//sample 305
i_data_q[49] = 9'd41;
i_data_i[50] = 9'd11;		//sample 306
i_data_q[50] =-9'd124;
i_data_i[51] = 9'd136;		//sample 307
i_data_q[51] = 9'd6;
i_data_i[52] = 9'd68;		//sample 308
i_data_q[52] = 9'd71;
i_data_i[53] = 9'd3;		//sample 309
i_data_q[53] =-9'd42;
i_data_i[54] =-9'd37;		//sample 310
i_data_q[54] = 9'd134;
i_data_i[55] =-9'd54;		//sample 311
i_data_q[55] =-9'd73;
i_data_i[56] =-9'd41;		//sample 312
i_data_q[56] =-9'd51;
i_data_i[57] =-9'd93;		//sample 313
i_data_q[57] =-9'd112;
i_data_i[58] =-9'd59;		//sample 314
i_data_q[58] =-9'd124;
i_data_i[59] =-9'd39;		//sample 315
i_data_q[59] = 9'd41;
i_data_i[60] = 9'd64;		//sample 316
i_data_q[60] = 9'd77;
i_data_i[61] = 9'd67;		//sample 317
i_data_q[61] = 9'd67;
i_data_i[62] = 9'd157;		//sample 318
i_data_q[62] =-9'd8;
i_data_i[63] =-9'd29;		//sample 319
i_data_q[63] = 9'd136;
#2
i_data_i[0] =-9'd124;		//sample 320
i_data_q[0] =-9'd28;
i_data_i[1] = 9'd73;		//sample 321
i_data_q[1] =-9'd64;
i_data_i[2] = 9'd68;		//sample 322
i_data_q[2] = 9'd72;
i_data_i[3] = 9'd132;		//sample 323
i_data_q[3] = 9'd74;
i_data_i[4] =-9'd75;		//sample 324
i_data_q[4] = 9'd112;
i_data_i[5] =-9'd48;		//sample 325
i_data_q[5] = 9'd36;
i_data_i[6] =-9'd41;		//sample 326
i_data_q[6] = 9'd17;
i_data_i[7] = 9'd18;		//sample 327
i_data_q[7] =-9'd116;
i_data_i[8] = 9'd89;		//sample 328
i_data_q[8] = 9'd84;
i_data_i[9] =-9'd82;		//sample 329
i_data_q[9] =-9'd32;
i_data_i[10] = 9'd93;		//sample 330
i_data_q[10] = 9'd26;
i_data_i[11] = 9'd10;		//sample 331
i_data_q[11] = 9'd157;
i_data_i[12] =-9'd68;		//sample 332
i_data_q[12] = 9'd1;
i_data_i[13] =-9'd34;		//sample 333
i_data_q[13] = 9'd156;
i_data_i[14] = 9'd15;		//sample 334
i_data_q[14] =-9'd65;
i_data_i[15] = 9'd23;		//sample 335
i_data_q[15] =-9'd36;
i_data_i[16] = 9'd60;		//sample 336
i_data_q[16] = 9'd85;
i_data_i[17] =-9'd37;		//sample 337
i_data_q[17] = 9'd118;
i_data_i[18] =-9'd46;		//sample 338
i_data_q[18] = 9'd87;
i_data_i[19] = 9'd77;		//sample 339
i_data_q[19] = 9'd100;
i_data_i[20] =-9'd58;		//sample 340
i_data_q[20] = 9'd61;
i_data_i[21] = 9'd79;		//sample 341
i_data_q[21] =-9'd70;
i_data_i[22] =-9'd67;		//sample 342
i_data_q[22] =-9'd104;
i_data_i[23] =-9'd41;		//sample 343
i_data_q[23] = 9'd95;
i_data_i[24] =-9'd3;		//sample 344
i_data_q[24] =-9'd132;
i_data_i[25] =-9'd72;		//sample 345
i_data_q[25] =-9'd41;
i_data_i[26] = 9'd3;		//sample 346
i_data_q[26] =-9'd104;
i_data_i[27] =-9'd91;		//sample 347
i_data_q[27] = 9'd14;
i_data_i[28] = 9'd51;		//sample 348
i_data_q[28] = 9'd80;
i_data_i[29] = 9'd51;		//sample 349
i_data_q[29] = 9'd40;
i_data_i[30] =-9'd92;		//sample 350
i_data_q[30] =-9'd39;
i_data_i[31] = 9'd100;		//sample 351
i_data_q[31] =-9'd88;
i_data_i[32] = 9'd20;		//sample 352
i_data_q[32] = 9'd42;
i_data_i[33] =-9'd121;		//sample 353
i_data_q[33] = 9'd35;
i_data_i[34] = 9'd77;		//sample 354
i_data_q[34] =-9'd57;
i_data_i[35] = 9'd84;		//sample 355
i_data_q[35] = 9'd15;
i_data_i[36] = 9'd137;		//sample 356
i_data_q[36] =-9'd1;
i_data_i[37] =-9'd17;		//sample 357
i_data_q[37] = 9'd129;
i_data_i[38] = 9'd39;		//sample 358
i_data_q[38] = 9'd84;
i_data_i[39] =-9'd114;		//sample 359
i_data_q[39] =-9'd39;
i_data_i[40] =-9'd54;		//sample 360
i_data_q[40] =-9'd19;
i_data_i[41] =-9'd85;		//sample 361
i_data_q[41] = 9'd37;
i_data_i[42] = 9'd103;		//sample 362
i_data_q[42] = 9'd107;
i_data_i[43] = 9'd37;		//sample 363
i_data_q[43] = 9'd15;
i_data_i[44] = 9'd90;		//sample 364
i_data_q[44] = 9'd61;
i_data_i[45] =-9'd50;		//sample 365
i_data_q[45] = 9'd102;
i_data_i[46] = 9'd61;		//sample 366
i_data_q[46] = 9'd87;
i_data_i[47] =-9'd133;		//sample 367
i_data_q[47] = 9'd14;
i_data_i[48] =-9'd8;		//sample 368
i_data_q[48] =-9'd117;
i_data_i[49] =-9'd14;		//sample 369
i_data_q[49] =-9'd47;
i_data_i[50] = 9'd137;		//sample 370
i_data_q[50] = 9'd34;
i_data_i[51] =-9'd5;		//sample 371
i_data_q[51] = 9'd98;
i_data_i[52] = 9'd25;		//sample 372
i_data_q[52] = 9'd93;
i_data_i[53] =-9'd47;		//sample 373
i_data_q[53] =-9'd12;
i_data_i[54] =-9'd25;		//sample 374
i_data_q[54] =-9'd76;
i_data_i[55] = 9'd113;		//sample 375
i_data_q[55] = 9'd96;
i_data_i[56] = 9'd49;		//sample 376
i_data_q[56] =-9'd93;
i_data_i[57] = 9'd89;		//sample 377
i_data_q[57] = 9'd67;
i_data_i[58] =-9'd107;		//sample 378
i_data_q[58] = 9'd41;
i_data_i[59] = 9'd112;		//sample 379
i_data_q[59] =-9'd33;
i_data_i[60] =-9'd37;		//sample 380
i_data_q[60] =-9'd144;
i_data_i[61] = 9'd34;		//sample 381
i_data_q[61] = 9'd89;
i_data_i[62] =-9'd51;		//sample 382
i_data_q[62] = 9'd8;
i_data_i[63] =-9'd66;		//sample 383
i_data_q[63] = 9'd87;
#2
i_data_i[0] =-9'd83;		//sample 384
i_data_q[0] = 9'd8;
i_data_i[1] =-9'd41;		//sample 385
i_data_q[1] =-9'd88;
i_data_i[2] = 9'd96;		//sample 386
i_data_q[2] =-9'd58;
i_data_i[3] = 9'd74;		//sample 387
i_data_q[3] =-9'd105;
i_data_i[4] =-9'd13;		//sample 388
i_data_q[4] =-9'd78;
i_data_i[5] =-9'd57;		//sample 389
i_data_q[5] = 9'd107;
i_data_i[6] =-9'd8;		//sample 390
i_data_q[6] =-9'd57;
i_data_i[7] =-9'd13;		//sample 391
i_data_q[7] =-9'd33;
i_data_i[8] =-9'd9;		//sample 392
i_data_q[8] = 9'd114;
i_data_i[9] =-9'd68;		//sample 393
i_data_q[9] =-9'd89;
i_data_i[10] = 9'd94;		//sample 394
i_data_q[10] =-9'd58;
i_data_i[11] = 9'd97;		//sample 395
i_data_q[11] =-9'd28;
i_data_i[12] =-9'd17;		//sample 396
i_data_q[12] = 9'd59;
i_data_i[13] = 9'd44;		//sample 397
i_data_q[13] = 9'd9;
i_data_i[14] =-9'd117;		//sample 398
i_data_q[14] =-9'd77;
i_data_i[15] = 9'd122;		//sample 399
i_data_q[15] = 9'd84;
i_data_i[16] =-9'd110;		//sample 400
i_data_q[16] = 9'd51;
i_data_i[17] = 9'd79;		//sample 401
i_data_q[17] = 9'd103;
i_data_i[18] =-9'd67;		//sample 402
i_data_q[18] = 9'd82;
i_data_i[19] =-9'd6;		//sample 403
i_data_q[19] = 9'd105;
i_data_i[20] =-9'd9;		//sample 404
i_data_q[20] = 9'd81;
i_data_i[21] = 9'd54;		//sample 405
i_data_q[21] =-9'd12;
i_data_i[22] =-9'd0;		//sample 406
i_data_q[22] =-9'd158;
i_data_i[23] = 9'd5;		//sample 407
i_data_q[23] =-9'd72;
i_data_i[24] =-9'd73;		//sample 408
i_data_q[24] = 9'd87;
i_data_i[25] = 9'd21;		//sample 409
i_data_q[25] =-9'd37;
i_data_i[26] = 9'd1;		//sample 410
i_data_q[26] =-9'd39;
i_data_i[27] =-9'd1;		//sample 411
i_data_q[27] =-9'd96;
i_data_i[28] = 9'd92;		//sample 412
i_data_q[28] = 9'd81;
i_data_i[29] =-9'd25;		//sample 413
i_data_q[29] = 9'd105;
i_data_i[30] = 9'd69;		//sample 414
i_data_q[30] = 9'd66;
i_data_i[31] =-9'd106;		//sample 415
i_data_q[31] = 9'd3;
i_data_i[32] = 9'd28;		//sample 416
i_data_q[32] =-9'd88;
i_data_i[33] =-9'd151;		//sample 417
i_data_q[33] = 9'd37;
i_data_i[34] = 9'd9;		//sample 418
i_data_q[34] = 9'd140;
i_data_i[35] = 9'd8;		//sample 419
i_data_q[35] =-9'd42;
i_data_i[36] =-9'd141;		//sample 420
i_data_q[36] =-9'd36;
i_data_i[37] =-9'd27;		//sample 421
i_data_q[37] = 9'd59;
i_data_i[38] =-9'd37;		//sample 422
i_data_q[38] = 9'd130;
i_data_i[39] =-9'd23;		//sample 423
i_data_q[39] = 9'd111;
i_data_i[40] =-9'd9;		//sample 424
i_data_q[40] = 9'd21;
i_data_i[41] =-9'd83;		//sample 425
i_data_q[41] = 9'd108;
i_data_i[42] = 9'd29;		//sample 426
i_data_q[42] =-9'd33;
i_data_i[43] = 9'd1;		//sample 427
i_data_q[43] = 9'd101;
i_data_i[44] = 9'd26;		//sample 428
i_data_q[44] =-9'd13;
i_data_i[45] = 9'd43;		//sample 429
i_data_q[45] = 9'd112;
i_data_i[46] = 9'd78;		//sample 430
i_data_q[46] = 9'd84;
i_data_i[47] = 9'd41;		//sample 431
i_data_q[47] = 9'd98;
i_data_i[48] =-9'd78;		//sample 432
i_data_q[48] = 9'd86;
i_data_i[49] =-9'd57;		//sample 433
i_data_q[49] =-9'd67;
i_data_i[50] = 9'd12;		//sample 434
i_data_q[50] = 9'd117;
i_data_i[51] =-9'd69;		//sample 435
i_data_q[51] = 9'd141;
i_data_i[52] = 9'd60;		//sample 436
i_data_q[52] =-9'd109;
i_data_i[53] = 9'd29;		//sample 437
i_data_q[53] =-9'd53;
i_data_i[54] = 9'd54;		//sample 438
i_data_q[54] =-9'd48;
i_data_i[55] = 9'd17;		//sample 439
i_data_q[55] = 9'd98;
i_data_i[56] = 9'd44;		//sample 440
i_data_q[56] =-9'd37;
i_data_i[57] =-9'd43;		//sample 441
i_data_q[57] = 9'd15;
i_data_i[58] =-9'd73;		//sample 442
i_data_q[58] =-9'd65;
i_data_i[59] =-9'd14;		//sample 443
i_data_q[59] =-9'd161;
i_data_i[60] = 9'd98;		//sample 444
i_data_q[60] =-9'd40;
i_data_i[61] = 9'd87;		//sample 445
i_data_q[61] =-9'd13;
i_data_i[62] = 9'd104;		//sample 446
i_data_q[62] =-9'd33;
i_data_i[63] =-9'd13;		//sample 447
i_data_q[63] =-9'd103;
#2
i_data_i[0] =-9'd11;		//sample 448
i_data_q[0] = 9'd119;
i_data_i[1] =-9'd20;		//sample 449
i_data_q[1] = 9'd101;
i_data_i[2] =-9'd98;		//sample 450
i_data_q[2] = 9'd27;
i_data_i[3] =-9'd4;		//sample 451
i_data_q[3] = 9'd117;
i_data_i[4] =-9'd33;		//sample 452
i_data_q[4] = 9'd7;
i_data_i[5] = 9'd46;		//sample 453
i_data_q[5] =-9'd2;
i_data_i[6] = 9'd118;		//sample 454
i_data_q[6] = 9'd8;
i_data_i[7] =-9'd70;		//sample 455
i_data_q[7] = 9'd56;
i_data_i[8] = 9'd85;		//sample 456
i_data_q[8] =-9'd58;
i_data_i[9] =-9'd21;		//sample 457
i_data_q[9] = 9'd41;
i_data_i[10] =-9'd46;		//sample 458
i_data_q[10] = 9'd120;
i_data_i[11] = 9'd42;		//sample 459
i_data_q[11] =-9'd116;
i_data_i[12] =-9'd22;		//sample 460
i_data_q[12] = 9'd41;
i_data_i[13] =-9'd108;		//sample 461
i_data_q[13] =-9'd6;
i_data_i[14] = 9'd41;		//sample 462
i_data_q[14] = 9'd103;
i_data_i[15] = 9'd86;		//sample 463
i_data_q[15] = 9'd55;
i_data_i[16] = 9'd32;		//sample 464
i_data_q[16] = 9'd96;
i_data_i[17] =-9'd12;		//sample 465
i_data_q[17] = 9'd103;
i_data_i[18] = 9'd1;		//sample 466
i_data_q[18] = 9'd39;
i_data_i[19] = 9'd39;		//sample 467
i_data_q[19] = 9'd10;
i_data_i[20] = 9'd103;		//sample 468
i_data_q[20] = 9'd45;
i_data_i[21] =-9'd10;		//sample 469
i_data_q[21] =-9'd38;
i_data_i[22] = 9'd90;		//sample 470
i_data_q[22] = 9'd52;
i_data_i[23] =-9'd94;		//sample 471
i_data_q[23] =-9'd7;
i_data_i[24] = 9'd105;		//sample 472
i_data_q[24] = 9'd10;
i_data_i[25] = 9'd118;		//sample 473
i_data_q[25] = 9'd9;
i_data_i[26] = 9'd107;		//sample 474
i_data_q[26] =-9'd57;
i_data_i[27] = 9'd29;		//sample 475
i_data_q[27] =-9'd49;
i_data_i[28] =-9'd97;		//sample 476
i_data_q[28] =-9'd63;
i_data_i[29] =-9'd5;		//sample 477
i_data_q[29] = 9'd87;
i_data_i[30] = 9'd72;		//sample 478
i_data_q[30] = 9'd45;
i_data_i[31] = 9'd58;		//sample 479
i_data_q[31] =-9'd24;
i_data_i[32] =-9'd121;		//sample 480
i_data_q[32] = 9'd26;
i_data_i[33] = 9'd36;		//sample 481
i_data_q[33] =-9'd106;
i_data_i[34] =-9'd138;		//sample 482
i_data_q[34] =-9'd8;
i_data_i[35] = 9'd27;		//sample 483
i_data_q[35] = 9'd106;
i_data_i[36] =-9'd64;		//sample 484
i_data_q[36] =-9'd27;
i_data_i[37] =-9'd110;		//sample 485
i_data_q[37] = 9'd6;
i_data_i[38] = 9'd88;		//sample 486
i_data_q[38] =-9'd131;
i_data_i[39] =-9'd115;		//sample 487
i_data_q[39] =-9'd97;
i_data_i[40] = 9'd102;		//sample 488
i_data_q[40] =-9'd29;
i_data_i[41] =-9'd80;		//sample 489
i_data_q[41] =-9'd135;
i_data_i[42] = 9'd64;		//sample 490
i_data_q[42] = 9'd70;
i_data_i[43] =-9'd67;		//sample 491
i_data_q[43] = 9'd97;
i_data_i[44] = 9'd62;		//sample 492
i_data_q[44] =-9'd68;
i_data_i[45] = 9'd41;		//sample 493
i_data_q[45] = 9'd101;
i_data_i[46] =-9'd83;		//sample 494
i_data_q[46] =-9'd44;
i_data_i[47] =-9'd94;		//sample 495
i_data_q[47] =-9'd70;
i_data_i[48] = 9'd38;		//sample 496
i_data_q[48] =-9'd130;
i_data_i[49] = 9'd115;		//sample 497
i_data_q[49] =-9'd6;
i_data_i[50] = 9'd52;		//sample 498
i_data_q[50] = 9'd17;
i_data_i[51] =-9'd46;		//sample 499
i_data_q[51] =-9'd37;
i_data_i[52] = 9'd105;		//sample 500
i_data_q[52] = 9'd51;
i_data_i[53] =-9'd93;		//sample 501
i_data_q[53] =-9'd128;
i_data_i[54] =-9'd12;		//sample 502
i_data_q[54] = 9'd107;
i_data_i[55] = 9'd2;		//sample 503
i_data_q[55] = 9'd116;
i_data_i[56] = 9'd60;		//sample 504
i_data_q[56] = 9'd60;
i_data_i[57] = 9'd37;		//sample 505
i_data_q[57] = 9'd7;
i_data_i[58] = 9'd11;		//sample 506
i_data_q[58] =-9'd33;
i_data_i[59] = 9'd118;		//sample 507
i_data_q[59] = 9'd16;
i_data_i[60] = 9'd64;		//sample 508
i_data_q[60] = 9'd61;
i_data_i[61] =-9'd37;		//sample 509
i_data_q[61] = 9'd139;
i_data_i[62] = 9'd47;		//sample 510
i_data_q[62] =-9'd2;
i_data_i[63] = 9'd93;		//sample 511
i_data_q[63] =-9'd37;
#2*/
for (j=0; j<64; j=j+1) begin 
	i_data_i[j] = 9'd0;		
	i_data_q[j] = 9'd0;
end
#(2*7)
	i_data_i[63] = 9'd128;
#2
	i_valid = 0;
	#40
    
	
	$finish;
end	

endmodule
